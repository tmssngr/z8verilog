`default_nettype none

module Memory #(
    parameter addrBusWidth = 8
) (
    input  wire                      clk,
    input  wire [addrBusWidth - 1:0] addr,
    input  wire                [7:0] dataIn,
    output reg                 [7:0] dataOut,
    input  wire                      write,
    input  wire                      strobe
);
    localparam size = 1 << addrBusWidth;
    reg [7:0] memory[0 : size - 1];
`ifdef BENCH
    integer i, file;
    initial begin
        for (i = 0; i < size; i = i + 1) begin
            memory[i] = 8'h0;
        end

        file = $fopen("memory.txt", "w");
    end
`endif

`include "alu.vh"
`include "assembly.vh"
`include "program.vh"
`ifdef BENCH
    initial begin
        $fclose(file);
    end
`endif
`include "sfr.vh"

    always @(posedge clk) begin
        if (strobe) begin
            if (write) begin
                memory[addr] <= dataIn;
                dataOut <= dataIn;
            end
            else begin
                dataOut <= memory[addr];
            end
        end
    end
endmodule

`include "Alu.v"

module Processor(
    input  wire        clk,
    //input  wire        reset,
    output wire [15:0] memAddr,
    input  wire  [7:0] memDataRead,
    output wire  [7:0] memDataWrite,
    output wire        memWrite,
    output wire        memStrobe,
    output wire  [7:0] port2Out,
    output wire  [3:0] port3Out
);
    `include "flags.vh"

    reg [15:0] pc, sp, addr;
    initial begin
        pc = 'hC;
        sp = 0;
    end

    reg  [7:0] instruction;
    wire [3:0] instrH = instruction[7:4];
    wire [3:0] instrL = instruction[3:0];
    wire isJumpRel = instrL == 4'hB;
    wire isJumpDA = instrL == 4'hD;
    wire isCallIRR = instrH == 4'hD && instrL == 4'h4;
    wire isCallDA = instrH == 4'hD && instrL == 4'h6;
    wire isInstrSize1 = instrL[3:1] == 3'b111;
    wire isInstrSize3 = ( (instrL[3:2] == 2'b01) // columns 04-07
                         | isJumpDA
                        ) & ~isCallIRR;
    wire isInstrSize2 = ~isInstrSize1 & ~isInstrSize3;

    reg  [7:0] second;
    wire [3:0] secondH = second[7:4];
    wire [3:0] secondL = second[3:0];

    reg  [7:0] third;
    wire [3:0] thirdH = third[7:4];
    wire [3:0] thirdL = third[3:0];
    wire [15:0] directAddress = {second, third};

    reg [3:0] rp = 0;
    reg [7:0] registers[0:'h7F];
    reg [7:0] p01m = 8'b01_0_01_1_01;
    //                  || | || | ++ P00-P03 Mode: 00 output, 01 input, 1x address A8-A11
    //                  || | || +--- Stack: 0 external,  1 internal
    //                  || | ++----- P1 Mode: 00 Output, 01 Input, 10 AD0-AD7, 11 tristate
    //                  || +-------- Memory timing: 0 normal, 1 extended
    //                  ++---------- P04-P07 Mode: 00 output, 01 input, 1x A12-A15 
    reg [7:0] p3m = 0;
    wire stackInternal = p01m[2];
    reg [7:0] port2;
    assign port2Out = port2;
    reg [7:0] port3;
    assign port3Out = port3[7:4];
    initial begin
        port2 = 0;
        port3 = 0;
        registers[2] = 0;
        registers[3] = 0;
    end

    reg [7:0] register;
    reg writeRegister = 0;

    `include "sfr.vh"
    `include "alu.vh"
    reg  [7:0] aluA = 0;
    reg  [7:0] aluB = 0;
    reg  [4:0] aluMode;
    wire [7:0] aluOut;
    reg  [7:0] flags = 0;
    wire [7:0] flagsOut;
    reg writeFlags = 0;
    Alu alu(
        .mode(aluMode),
        .a(aluA),
        .b(aluB),
        .flags(flags),
        .out(aluOut),
        .outFlags(flagsOut)
    );

    function [7:0] r4(
        input [3:0] r
    );
        r4 = { rp, r };
    endfunction

    function [7:0] r8(
        input [7:0] r
    );
        if (r[7:4] == 4'hE)
            r8 = r4(r[3:0]);
        else
            r8 = r;
    endfunction

    function [7:0] readRegister8(
        input [7:0] r
    );
        casez (r)
        2:            readRegister8 = port2;
        3:            readRegister8 = port3;
        8'b0???_????: readRegister8 = registers[r[6:0]];
        P01M:         readRegister8 = p01m;
        P3M:          readRegister8 = p3m;
        FLAGS:        readRegister8 = flags;
        RP:           readRegister8 = { rp, 4'h0 };
        SPH:          readRegister8 = sp[15:8];
        SPL:          readRegister8 = sp[7:0];
        default:      readRegister8 = 0;
        endcase
    endfunction

    function [7:0] readRegister4(
        input [3:0] r
    );
        readRegister4 = readRegister8(r4(r));
    endfunction

    function [4:0] alu1OpCode(
        input[3:0] instrH
    );
        alu1OpCode = { 1'b0, instrH };
    endfunction

    function [4:0] alu2OpCode(
        input[3:0] instrH
    );
        alu2OpCode = { 1'b1, instrH };
    endfunction

    reg takeBranchTmp;
    always @(*) begin
        case (instrH[2:0])
        0: takeBranchTmp = 0;
        1: takeBranchTmp =  flags[FLAG_INDEX_S] ^ flags[FLAG_INDEX_V];
        2: takeBranchTmp = (flags[FLAG_INDEX_S] ^ flags[FLAG_INDEX_V]) | flags[FLAG_INDEX_Z];
        3: takeBranchTmp =  flags[FLAG_INDEX_C] | flags[FLAG_INDEX_Z];
        4: takeBranchTmp =  flags[FLAG_INDEX_V];
        5: takeBranchTmp =  flags[FLAG_INDEX_S];
        6: takeBranchTmp =  flags[FLAG_INDEX_Z];
        7: takeBranchTmp =  flags[FLAG_INDEX_C];
        endcase
    end
    wire takeBranch = takeBranchTmp ^ instrH[3];

`ifdef BENCH
    function [1:4*8] alu1OpName(
        input [3:0] instrH
    );
    begin
        case (instrH)
        ALU1_DEC : alu1OpName = "dec";
        ALU1_RLC : alu1OpName = "rlc";
        ALU1_INC : alu1OpName = "inc";
        ALU1_DA  : alu1OpName = "da";
        ALU1_COM : alu1OpName = "com";
        ALU1_DECW: alu1OpName = "decw";
        ALU1_RL  : alu1OpName = "rl";
        ALU1_INCW: alu1OpName = "incw";
        ALU1_CLR : alu1OpName = "clr";
        ALU1_RRC : alu1OpName = "rrc";
        ALU1_SRA : alu1OpName = "sra";
        ALU1_RR  : alu1OpName = "rr";
        ALU1_SWAP: alu1OpName = "swap";
        default  : alu1OpName = "?";
        endcase;
    end
    endfunction

    function [1:3*8] alu2OpName(
        input [3:0] instrH
    );
    begin
        case (alu2OpCode(instrH))
        ALU2_ADD: alu2OpName = "add";
        ALU2_ADC: alu2OpName = "adc";
        ALU2_SUB: alu2OpName = "sub";
        ALU2_SBC: alu2OpName = "sbc";
        ALU2_OR : alu2OpName = "or";
        ALU2_AND: alu2OpName = "and";
        ALU2_TCM: alu2OpName = "tcm";
        ALU2_TM : alu2OpName = "tm";
        ALU2_CP : alu2OpName = "cp";
        ALU2_XOR: alu2OpName = "xor";
        default : alu2OpName = "?";
        endcase
    end
    endfunction

    function [1:3*8] ccName(
        input [3:0] instrH
    );
    begin
        case (instrH)
        0: ccName = "f";
        1: ccName = "lt";
        2: ccName = "le";
        3: ccName = "ule";
        4: ccName = "ov";
        5: ccName = "mi";
        6: ccName = "z";
        7: ccName = "c";
        8: ccName = "";
        9: ccName = "ge";
        10: ccName = "gt";
        11: ccName = "ugt";
        12: ccName = "nov";
        13: ccName = "pl";
        14: ccName = "nz";
        15: ccName = "nc";
        endcase
    end
    endfunction
`endif

    `include "states.vh"
    reg [FETCH_MSB:0] fetchState = FETCH_INSTR_WAIT;
    reg [OP_MSB:0] opType = OP_UNDECIDED;
    reg [OPSTATE_MSB:0] opState = OPSTATE0;

    wire [15:0] nextRelativePc = pc + { {8{second[7]}}, second };
    wire [15:0] nextPc = ( fetchState == FETCH_INSTR_READ
                         | fetchState == FETCH_SECOND_READ
                         | fetchState == FETCH_THIRD_READ
                         ) ? pc + 16'b1
                           : ( (fetchState == FETCH_DECODE & isJumpRel & takeBranch)
                             || (opType == OP_DJNZ & opState == OPSTATE2)
                             ) ? nextRelativePc
                               : ( (opType == OP_RET  & opState == OPSTATE5)
                                 | (opType == OP_CALL & opState == OPSTATE6)
                                 | (opType == OP_JP   & opState == OPSTATE2)
                                 ) ? addr
                                   : pc;
    reg readMem = 0;
    reg writeMem = 0;
    assign memAddr = readMem | writeMem
                     ? addr : pc;
    assign memDataWrite = aluA;
    assign memWrite = writeMem;
    assign memStrobe = (fetchState == FETCH_INSTR_WAIT)
                     | (fetchState == FETCH_SECOND_WAIT & ~isInstrSize1)
                     | (fetchState == FETCH_THIRD_WAIT)
                     | readMem
                     | writeMem;
`ifdef BENCH
    reg[4:0] cycleCounter = 0;
    reg[4:0] expectedCycles = 0;
`endif

    task nextCommand;
        begin
            fetchState <= FETCH_INSTR_WAIT;
            opState <= OPSTATE0;
            opType <= OP_UNDECIDED;
        end
    endtask

    always @(posedge clk) begin
        if (writeFlags) begin
`ifdef BENCH
            $display("    alu:    %h       %h    =>    %h", aluA, aluB, aluOut);
            $display("         %b %b => %b", aluA, aluB, aluOut);
            $display("    flags = %b_%b", flagsOut[7:4], flagsOut[3:0]);
`endif
            flags <= flagsOut;
        end
        writeFlags <= 0;

        if (writeRegister) begin
`ifdef BENCH
            $display("    reg[%h] = %h", register, aluOut);
`endif
            casez (register)
            8'b0???_????: registers[register] <= aluOut;
            P01M:         p01m                <= aluOut;
            P3M:          p3m                 <= aluOut;
            FLAGS:        flags               <= aluOut;
            RP:           rp                  <= aluOut[7:4];
            SPH:          sp[15:8]            <= aluOut;
            SPL:          sp[7:0]             <= aluOut;
            endcase

            // store in registers AND ports, so it is easier to check registers
            case (register)
            2: port2 <= aluOut;
            3: port3 <= aluOut;
            endcase
        end
        writeRegister <= 0;
        readMem <= 0;
        writeMem <= 0;

`ifdef BENCH
        if (fetchState == FETCH_INSTR_WAIT) begin
            if (cycleCounter != 0) begin
                if (expectedCycles == 0) begin
                    $display("expected cycles not defined");
                    $finish(2);
                end

                if (cycleCounter < expectedCycles) 
                    $display("%d cycles, expected %d", cycleCounter, expectedCycles);
                else if (cycleCounter > expectedCycles) 
                    $display("%d cycles, expected %d - TOO SLOW", cycleCounter, expectedCycles);
                else
                    $display("exact %d cycles", cycleCounter);
                expectedCycles <= 0;
            end
            cycleCounter <= 1;
        end
        else begin
            cycleCounter <= cycleCounter + 1;
        end
`endif

        if (fetchState != FETCH_DECODE) begin
            fetchState <= fetchState + FETCH_INC;
        end
        if (opType != OP_UNDECIDED) begin
            opState <= opState + OPSTATE_INC;
        end

        case (fetchState)
        FETCH_INSTR_WAIT: begin
`ifdef BENCH
            addr <= 0;
            aluA <= 0;
            aluB <= 0;
            aluMode <= 0;
            register <= 0;
            instruction <= 0;
            second <= 0;
            third <= 0;
`endif
        end

        FETCH_INSTR_READ: begin
`ifdef BENCH
            $display("\n%h: read 1st byte %h", pc, memDataRead);
`endif
            instruction <= memDataRead;
        end

        FETCH_SECOND_WAIT: begin
            if (isInstrSize1) begin
                fetchState <= FETCH_DECODE;
            end
        end

        FETCH_SECOND_READ: begin
`ifdef BENCH
            $display("%h: read 2nd byte %h", pc, memDataRead);
`endif
            second <= memDataRead;
            if (isInstrSize2) begin
                fetchState <= FETCH_DECODE;
            end
        end

        FETCH_THIRD_WAIT: begin
        end

        FETCH_THIRD_READ: begin
`ifdef BENCH
            $display("%h: read 3rd byte %h", pc, memDataRead);
`endif
            third <= memDataRead;
        end

        FETCH_DECODE: begin
            if (opType == OP_UNDECIDED) begin
    `ifdef BENCH
                // $display("  decoding");
                if (isInstrSize1)
                    $display("  %h", instruction);
                else if (isInstrSize2)
                    $display("  %h %h", instruction, second);
                else if (isInstrSize3)
                    $display("  %h %h %h", instruction, second, third);
    `endif
                case (instrL)
                // ================================================================
                // Column 0
                // ================================================================
                4'h0: begin
                    case (instrH)
                    4'h3: begin
    `ifdef BENCH
                        $display("    jp @%h", second);
                        expectedCycles <= 8;
    `endif
                        opType <= OP_JP;
                    end
                    4'h5: begin
    `ifdef BENCH
                        $display("    pop %h", second);
                        expectedCycles <= 10;
    `endif
                        // dst <- @SP
                        // SP <- SP + 1
                        register <= r8(second);
                        opType <= OP_POP;
                    end
                    4'h7: begin
    `ifdef BENCH
                        $display("    push %h", second);
                        expectedCycles <= stackInternal ? 10 : 12;
    `endif
                        register <= r8(second);
                        opType <= stackInternal 
                            ? OP_PUSH_I
                            : OP_PUSH_E;
                    end
                    4'h8: begin
    `ifdef BENCH
                        $display("    decw %h", second);
                        expectedCycles <= 10;
    `endif
                        opType <= OP_ALU1WORD;
                    end
                    4'hA: begin
    `ifdef BENCH
                        $display("    incw %h", second);
                        expectedCycles <= 10;
    `endif
                        opType <= OP_ALU1WORD;
                    end
                    default: begin
    `ifdef BENCH
                        $display("   %s %h", 
                                alu1OpName(instrH), second);
                        expectedCycles <= instrH == 4 ? 8 : 6;
    `endif
                        aluMode <= alu1OpCode(instrH);
                        register <= r8(second);
                        opType <= OP_ALU1;
                    end
                    endcase
                end
                // ================================================================
                // Column 1
                // ================================================================
                4'h1: begin
                    case (instrH)
                    4'h3: begin
    `ifdef BENCH
                        $display("    srp %h", second);
                        expectedCycles <= 6;
    `endif
                        register <= RP;
                        opType <= OP_LD;
                    end
                    4'h5: begin
    `ifdef BENCH
                        $display("    pop @%h", second);
                        expectedCycles <= 10;
    `endif
                        register <= readRegister8(r8(second));
                        opType <= OP_POP;
                    end
                    4'h7: begin
    `ifdef BENCH
                        $display("    push @%h", second);
                        expectedCycles <= stackInternal ? 12 : 14;
    `endif
                        register <= readRegister8(r8(second));
                        opType <= stackInternal 
                            ? OP_PUSH_I
                            : OP_PUSH_E;
                    end
                    4'h8: begin
    `ifdef BENCH
                        $display("    decw @%h", second);
                        expectedCycles <= 10;
    `endif
                        opType <= OP_ALU1WORD;
                    end
                    4'hA: begin
    `ifdef BENCH
                        $display("    incw @%h", second);
                        expectedCycles <= 10;
    `endif
                        opType <= OP_ALU1WORD;
                    end
                    default: begin
    `ifdef BENCH
                        $display("   %s @%h", 
                                alu1OpName(instrH), second);
                        expectedCycles <= instrH == 4 ? 8 : 6;
    `endif
                        aluMode <= alu1OpCode(instrH);
                        register <= readRegister8(r8(second));
                        opType <= OP_ALU1;
                    end
                    endcase
                end
                // ================================================================
                // Column 2
                // ================================================================
                4'h2: begin
                    case (instrH)
                    4'h8: begin
    `ifdef BENCH
                        $display("    lde r%h, Irr%h",
                                secondH, secondL);
                        expectedCycles <= 12;
    `endif
                        register <= r4(secondH);
                        opType <= OP_LDC;
                    end
                    4'h9: begin
    `ifdef BENCH
                        $display("    lde Irr%h, r%h",
                                secondL, secondH);
                        expectedCycles <= 12;
    `endif
                        register <= r4(secondH);
                        opType <= OP_LDC;
                    end
                    4'hC: begin
    `ifdef BENCH
                        $display("    ldc r%h, Irr%h",
                                secondH, secondL);
                        expectedCycles <= 12;
    `endif
                        register <= r4(secondH);
                        opType <= OP_LDC;
                    end
                    4'hD: begin
    `ifdef BENCH
                        $display("    ldc Irr%h, r%h",
                                secondL, secondH);
                        expectedCycles <= 12;
    `endif
                        register <= r4(secondH);
                        opType <= OP_LDC;
                    end
                    4'hE,
                    4'hF: begin
    `ifdef BENCH
                        $display("    ? %h", second);
    `endif
                        opType <= OP_ILLEGAL;
                    end
                    // x2
                    default: begin
    `ifdef BENCH
                        $display("    %s r%h, r%h",
                                alu2OpName(instrH),
                                secondH, secondL);
                        expectedCycles <= 6;
    `endif
                        register <= r4(secondL);
                        opType <= OP_ALU2;
                    end
                    endcase
                end
                // ================================================================
                // Column 3
                // ================================================================
                4'h3: begin
                    case (instrH)
                    4'h8: begin
    `ifdef BENCH
                        $display("    ldei Ir%h, Irr%h",
                                secondH, secondL);
                        expectedCycles <= 18;
    `endif
                        register <= readRegister4(secondH);
                        opType <= OP_LDC;
                    end
                    4'h9: begin
    `ifdef BENCH
                        $display("    ldei Irr%h, Ir%h",
                                secondL, secondH);
                        expectedCycles <= 18;
    `endif
                        register <= readRegister4(secondH);
                        opType <= OP_LDC;
                    end
                    4'hC: begin
    `ifdef BENCH
                        $display("    ldci Ir%h, Irr%h",
                                secondH, secondL);
                        expectedCycles <= 18;
    `endif
                        register <= readRegister4(secondH);
                        opType <= OP_LDC;
                    end
                    4'hD: begin
    `ifdef BENCH
                        $display("    ldci Irr%h, Ir%h",
                                secondL, secondH);
                        expectedCycles <= 18;
    `endif
                        register <= readRegister4(secondH);
                        opType <= OP_LDC;
                    end
                    4'hE: begin
    `ifdef BENCH
                        $display("    ld r%h, @r%h",
                                secondH, secondL);
                        expectedCycles <= 6;
    `endif
                        register <= readRegister4(secondL);
                        opType <= OP_LD;
                    end
                    4'hF: begin
    `ifdef BENCH
                        $display("    ld @r%h, r%h",
                                secondH, secondL);
                        expectedCycles <= 6;
    `endif
                        register <= readRegister4(secondH);
                        opType <= OP_LD;
                    end
                    default: begin
    `ifdef BENCH
                        $display("    %s r%h, Ir%h",
                                alu2OpName(instrH),
                                secondH, secondL);
                        expectedCycles <= 6;
    `endif
                        register <= readRegister4(secondL);
                        opType <= OP_ALU2;
                    end
                    endcase
                end
                // ================================================================
                // Column 4
                // ================================================================
                4'h4: begin
                    case (instrH)
                    4'h8,
                    4'h9,
                    4'hC,
                    4'hF: begin
    `ifdef BENCH
                        $display("    ? %h", instruction);
    `endif
                        opType <= OP_ILLEGAL;
                    end
                    4'hD: begin
    `ifdef BENCH
                        $display("    call @%h", second);
                        expectedCycles <= 20;
    `endif
                        opType <= OP_CALL;
                    end
                    4'hE: begin
    `ifdef BENCH
                        $display("    ld %h, %h", third, second);
                        expectedCycles <= 10;
    `endif
                        register <= r8(second);
                        opType <= OP_LD;
                    end
                    // x4
                    default: begin
    `ifdef BENCH
                        $display("    %s %h, %h",
                                alu2OpName(instrH),
                                third, second);
                        expectedCycles <= 10;
    `endif
                        register <= r8(second);
                        opType <= OP_ALU2;
                    end
                    endcase
                end
                // ================================================================
                // Column 5
                // ================================================================
                4'h5: begin
                    case (instrH)
                    4'h8,
                    4'h9,
                    4'hC,
                    4'hD:
                    begin
    `ifdef BENCH
                        $display("    ? %h", instruction);
    `endif
                        opType <= OP_ILLEGAL;
                    end
                    4'hE: begin
    `ifdef BENCH
                        $display("    ld %h, @%h", third, second);
                        expectedCycles <= 10;
    `endif
                        register <= readRegister8(r8(second));
                        opType <= OP_LD;
                    end
                    4'hF: begin
    `ifdef BENCH
                        $display("    ld @%h, %h", third, second);
                        expectedCycles <= 10;
    `endif
                        aluA <= readRegister8(r8(second));
                        opType <= OP_LD;
                    end
                    // x5
                    default: begin
    `ifdef BENCH
                        $display("    %s %h, @%h",
                                alu2OpName(instrH),
                                third, second);
                        expectedCycles <= 10;
    `endif
                        register <= readRegister8(r8(second));
                        opType <= OP_ALU2;
                    end
                    endcase
                end
                // ================================================================
                // Column 6
                // ================================================================
                4'h6: begin
                    case (instrH)
                    4'h8,
                    4'h9,
                    4'hC,
                    4'hF: begin
    `ifdef BENCH
                        $display("    ? %h", instruction);
    `endif
                        opType <= OP_ILLEGAL;
                    end
                    4'hD: begin
    `ifdef BENCH
                        $display("    call %h", directAddress);
                        expectedCycles <= 20;
    `endif
                        opType <= OP_CALL;
                    end
                    4'hE: begin
    `ifdef BENCH
                        $display("    ld %h, #%h", second, third);
                        expectedCycles <= 10;
    `endif
                        register <= r8(second);
                        opType <= OP_LD;
                    end
                    default: begin
    `ifdef BENCH
                        $display("    %s %h, #%h",
                                alu2OpName(instrH),
                                second, third);
                        expectedCycles <= 10;
    `endif
                        register <= r8(second);
                        opType <= OP_ALU2;
                    end
                    endcase
                end
                // ================================================================
                // Column 7
                // ================================================================
                4'h7: begin
                    case (instrH)
                    4'h8,
                    4'h9,
                    4'hF: begin
    `ifdef BENCH
                        $display("    ? %h", instruction);
    `endif
                        opType <= OP_ILLEGAL;
                    end
                    4'hC: begin
    `ifdef BENCH
                        $display("    ld r%h, @r%h+%h", 
                                secondH, secondL, third);
                        expectedCycles <= 10;
    `endif
                        register <= readRegister4(secondL);
                        opType <= OP_LD;
                    end
                    4'hD: begin
    `ifdef BENCH
                        $display("    ld @r%h+%h, r%h", 
                                secondL, third, secondH);
                        expectedCycles <= 10;
    `endif
                        register <= readRegister4(secondL);
                        opType <= OP_LD;
                    end
                    4'hE: begin
    `ifdef BENCH
                        $display("    ld @%h, #%h", second, third);
                        expectedCycles <= 10;
    `endif
                        register <= readRegister8(r8(second));
                        opType <= OP_LD;
                    end
                    default: begin
    `ifdef BENCH
                        $display("    %s @%h, #%h",
                                alu2OpName(instrH),
                                second, third);
                        expectedCycles <= 10;
    `endif
                        register <= readRegister8(r8(second));
                        opType <= OP_ALU2;
                    end
                    endcase
                end
                // ================================================================
                // Column 8
                // ================================================================
                4'h8: begin
    `ifdef BENCH
                    $display("    ld r%h, %h", instrH, second);
                    expectedCycles <= 6;
    `endif
                    register <= r4(instrH);
                    opType <= OP_LD;
                end
                // ================================================================
                // Column 9
                // ================================================================
                4'h9: begin
    `ifdef BENCH
                    $display("    ld %h, r%h", second, instrH);
                    expectedCycles <= 6;
    `endif
                    register <= second; // no r8(second) !
                    opType <= OP_LD;
                end
                // ================================================================
                // Column A
                // ================================================================
                4'hA: begin
    `ifdef BENCH
                    $display("    djnz r%h, %h", instrH, second);
    `endif
                    register <= r4(instrH);
                    opType <= OP_DJNZ;
                end
                // ================================================================
                // Column B
                // ================================================================
                4'hB: begin
    `ifdef BENCH
                    $display("    jr %s, %h", ccName(instrH), second);
                    expectedCycles <= takeBranch ? 12 : 10;
    `endif
                    nextCommand();
                end
                // ================================================================
                // Column C
                // ================================================================
                4'hC: begin
    `ifdef BENCH
                    $display("    ld r%h, #%h", instrH, second);
                    expectedCycles <= 6;
    `endif
                    register <= r4(instrH);
                    opType <= OP_LD;
                end
                // ================================================================
                // Column D
                // ================================================================
                4'hD: begin
    `ifdef BENCH
                    $display("    jp %s, %h", ccName(instrH), directAddress);
                    expectedCycles <= takeBranch ? 12 : 10;
    `endif
                    if (takeBranch)
                        opType <= OP_JP;
                    else
                        nextCommand();
                end
                // ================================================================
                // Column E
                // ================================================================
                4'hE: begin
    `ifdef BENCH
                    $display("    inc r%h", instrH);
                    expectedCycles <= 6;
    `endif
                    register <= r4(instrH);
                    aluMode <= ALU1_INC;
                    opType <= OP_ALU1;
                end
                // ================================================================
                // Column F
                // ================================================================
                4'hF: begin
                    case (instrH)
                    4'h8: begin
    `ifdef BENCH
                        $display("    di");
                        expectedCycles <= 6;
    `endif
                        //TODO
                        nextCommand();
                    end
                    4'h9: begin
    `ifdef BENCH
                        $display("    ei");
                        expectedCycles <= 6;
    `endif
                        //TODO
                        nextCommand();
                    end
                    4'hA: begin
    `ifdef BENCH
                        $display("    ret");
                        expectedCycles <= 14;
    `endif
                        opType <= OP_RET;
                    end
                    4'hB: begin
    `ifdef BENCH
                        $display("    iret");
                        expectedCycles <= 16;
    `endif
                        opType <= OP_IRET;
                    end
                    4'hC: begin
    `ifdef BENCH
                        $display("    rcf");
                        expectedCycles <= 6;
    `endif
                        flags[FLAG_INDEX_C] <= instrH[0];
                        nextCommand();
                    end
                    4'hD: begin
    `ifdef BENCH
                        $display("    scf");
                        expectedCycles <= 6;
    `endif
                        flags[FLAG_INDEX_C] <= instrH[0];
                        nextCommand();
                    end
                    4'hE: begin
    `ifdef BENCH
                        $display("    ccf");
                        expectedCycles <= 6;
    `endif
                        flags[FLAG_INDEX_C] <= ~flags[FLAG_INDEX_C];
                        nextCommand();
                    end
                    4'hF: begin
    `ifdef BENCH
                        $display("    nop");
                        expectedCycles <= 6;
    `endif
                        nextCommand();
                    end
                    default: begin
    `ifdef BENCH
                        $display("    ?");
    `endif
                        opType <= OP_ILLEGAL;
                    end
                    endcase
                end
                default: begin
                end
                endcase
            end
        end
    endcase

    case (opType)
        OP_LD: begin
            case (instrL)
            4'h1: begin
                // srp
                aluA <= second;
            end
            4'h3: begin
                case (instrH)
                4'hE: begin
                    aluA <= readRegister8(register);
                    register <= r4(secondH);
                end
                4'hF: begin
                    aluA <= readRegister4(secondL);
                end
                endcase
            end
            4'h4: begin
                case (instrH)
                4'hE: begin
                    aluA <= readRegister8(register);
                    register <= r8(third);
                end
                endcase
            end
            4'h5: begin
                case (instrH)
                4'hE: begin
                    aluA <= readRegister8(register);
                    register <= r8(third);
                end
                4'hF: begin
                    register <= readRegister8(r8(third));
                end
                endcase
            end
            4'h6: begin
                case (instrH)
                4'hE: begin
                    aluA <= third;
                end
                endcase
            end
            4'h7: begin
                case (instrH)
                4'hC: begin
                    aluA <= readRegister8(register + third);
                    register <= r4(secondH);
                end
                4'hD: begin
                    aluA <= readRegister4(secondH);
                    register <= register + third;
                end
                4'hE: begin
                    aluA <= third;
                end
                endcase
            end
            4'h8: begin
                aluA <= readRegister8(r8(second));
            end
            4'h9: begin
                aluA <= readRegister4(instrH);
            end
            4'hC: begin
                aluA <= second;
            end
            endcase
            aluMode <= ALU1_LD;
            writeRegister <= 1;
            nextCommand();
        end
        OP_ALU1: begin
            case (opState)
            OPSTATE0: begin
                aluA <= readRegister8(register);
                writeRegister <= 1;
                writeFlags <= 1;

                if (aluMode != ALU1_DA)
                    nextCommand();
            end
            default: begin
                aluA <= aluOut;
                aluMode <= ALU1_DA_H;
                writeRegister <= 1;
                writeFlags <= 1;
                nextCommand();
            end
            endcase
        end
        OP_ALU1WORD: begin
            case (opState)
            OPSTATE0: begin
                aluMode <= instrH & 7;
                register <= instrL & 1 
                    ? readRegister8(r8(second))
                    : r8(second);
            end
            OPSTATE1: begin
                register <= {register[7:1], 1'h1};
            end
            OPSTATE2: begin
                aluA <= readRegister8(register);
                writeRegister <= 1;
            end
            OPSTATE3: begin
                register <= { register[7:1], 1'b0 };
            end
            default: begin
                aluA <= readRegister8(register);
                aluB <= aluOut;
                aluMode <= aluMode | 'h8; // inc/dec -> incw/decw
                writeRegister <= 1;
                writeFlags <= 1;
                nextCommand();
            end
            endcase
        end
        OP_ALU2: begin
            case (opState)
            OPSTATE0: begin
                case (instrL)
                2, // r, r
                3: // r, Ir
                begin
                    aluB <= readRegister8(register);
                    register <= r4(secondH);
                end
                4, // R, R
                5: // R, IR
                begin
                    aluB <= readRegister8(register);
                    register <= r8(third);
                end
                6, // R, IM
                7: // IR, IM
                begin
                    aluB <= third;
                end
                endcase
            end
            OPSTATE1: begin
                aluA <= readRegister8(register);
            end
            default: begin
                aluMode <= alu2OpCode(instrH);
                writeRegister <= (instrH[3:2] == 2'b00)     // add, adc, sub, sbc
                                | (instrH[3:1] == 3'b010)   // or, and
                                | (instrH      == 4'b1011); // xor
                writeFlags <= 1;
                nextCommand();
            end
            endcase
        end
        OP_POP: begin
            case (opState)
            OPSTATE0: begin
                addr <= sp;
                readMem <= 1;
            end
            OPSTATE1: begin
                readMem <= 1;
            end
            OPSTATE2: begin
                aluA <= stackInternal
                    ? readRegister8(addr[7:0])
                    : memDataRead;
            end
            default: begin
                aluMode <= ALU1_LD;
                sp <= sp + 16'b1;
                writeRegister <= 1;
                nextCommand();
            end
            endcase
        end
        OP_PUSH_I: begin
            case (opState)
            OPSTATE0: begin
                sp <= sp - 16'b1;
            end
            default: begin
                aluMode <= ALU1_LD;
                aluA <= readRegister8(register);
                register <= sp[7:0];
                writeRegister <= 1;
                nextCommand();
            end
            endcase
        end
        OP_PUSH_E: begin
            case (opState)
            OPSTATE0: begin
                sp <= sp - 16'b1;
            end
            OPSTATE1: begin
                aluA <= readRegister8(register);
                addr <= sp;
                writeMem <= 1;
            end
            default: begin
                nextCommand();
            end
            endcase
        end
        OP_DJNZ: begin
            case (opState)
            OPSTATE0: begin
                aluA <= readRegister8(register);
                aluMode <= ALU1_DEC;
                writeRegister <= 1;
            end
            OPSTATE1: begin
`ifdef BENCH
                expectedCycles <= flagsOut[FLAG_INDEX_Z] ? 10 : 12;
`endif
                if (flagsOut[FLAG_INDEX_Z])
                    nextCommand();
            end
            default: begin
                nextCommand();
            end
            endcase
        end
        OP_JP: begin
            case (opState)
            OPSTATE0: begin
                addr[15:8] = isJumpDA
                    ? second
                    : readRegister8(r8({second[7:1], 1'b0}));
            end
            OPSTATE1: begin
                addr[7:0] = isJumpDA
                    ? third
                    : readRegister8(r8({second[7:1], 1'b1}));
            end
            default: begin
                nextCommand();
            end
            endcase
        end
        OP_CALL: begin
            // push PCL, PCH
            case (opState)
            OPSTATE0: begin
                sp <= sp - 16'b1;
                aluA <= pc[7:0];
            end
            OPSTATE1,
            OPSTATE3: begin
                if (stackInternal) begin
                    aluMode <= ALU1_LD;
                    register <= sp[7:0];
                    writeRegister <= 1;
                end
                else begin
                    addr <= sp;
                    writeMem <= 1;
                end
            end
            OPSTATE2: begin
                sp <= sp - 16'b1;
                aluA <= pc[15:8];
            end
            OPSTATE4: begin
                addr[15:8] = isCallDA 
                    ? second
                    : readRegister8(r8({second[7:1], 1'b0}));
            end
            OPSTATE5: begin
                addr[7:0] = isCallDA
                    ? third
                    : readRegister8(r8({second[7:1], 1'b1}));
            end
            default: begin
                nextCommand();
            end
            endcase
        end
        OP_IRET: begin
            // flags, PCH, PCL
            case (opState)
            OPSTATE0: begin
                addr <= sp;
                sp <= sp + 16'b1;
                readMem <= ~stackInternal;
            end
            OPSTATE1: begin
                aluMode <= ALU1_LD;
                aluA <= stackInternal
                    ? readRegister8(addr[7:0])
                    : memDataRead;
                register <= FLAGS;
                writeRegister <= 1;
                opType <= OP_RET;
                opState <= OPSTATE0;
            end
            endcase
        end
        OP_RET: begin
            // PCH, PCL
            case (opState)
            OPSTATE0: begin
                addr <= sp;
                readMem <= ~stackInternal;
            end
            OPSTATE1: begin
                sp <= sp + 16'b1;
                readMem <= ~stackInternal;
            end
            OPSTATE2: begin
                aluA <= stackInternal
                    ? readRegister8(addr[7:0])
                    : memDataRead;// temp
                addr <= sp;
                readMem <= ~stackInternal;
            end
            OPSTATE3: begin
                sp <= sp + 16'b1;
                readMem <= ~stackInternal;
            end
            OPSTATE4: begin
                addr[15:8] <= aluA;
                addr[7:0] <= stackInternal
                    ? readRegister8(addr[7:0])
                    : memDataRead;
            end
            default: begin
                nextCommand();
                //TODO: for iret enable interrupts
            end
            endcase
        end
        OP_LDC: begin
            case (opState)
            OPSTATE0: begin
                addr[15:8] <= readRegister4({secondL[3:1], 1'b0});
            end
            OPSTATE1: begin
                addr[7:0] <= readRegister4({secondL[3:1], 1'b1});
                if (instrH[0] == 0)
                    readMem <= 1;
            end
            OPSTATE2: begin
                if (instrH[0] == 0) begin
                    readMem <= 1;
                end
                else begin
                    aluA <= readRegister8(register);
                    writeMem <= 1;
                end
            end
            OPSTATE3: begin
                if (instrH[0] == 0) begin
                    aluA <= memDataRead;
                    aluMode <= ALU1_LD;
                    writeRegister <= 1;
                end
                // ldci?
                if (instrL[0] == 0)
                    nextCommand();
            end
            OPSTATE4: begin
                aluA <= register;
                register <= r4(secondH);
                aluMode <= ALU1_INC;
                writeRegister <= 1;
            end
            OPSTATE5: begin
                aluA <= addr[7:0];
                register <= r4({secondL[3:1], 1'b1});
                aluMode <= ALU1_INC;
                writeRegister <= 1;
            end
            OPSTATE6: begin
                aluA <= addr[15:8];
                aluB <= aluOut;
                register[0] <= 1'b0;
                aluMode <= ALU1_INCW;
                writeRegister <= 1;
                nextCommand();
            end
            endcase
        end
        OP_ILLEGAL: begin
            opState <= OPSTATE0;
        end
        endcase
        pc <= nextPc;
    end
endmodule

module SoC(
    input  wire       clk,
    output wire [7:0] port2,
    output wire [3:0] port3
);
    wire [15:0] memAddr;
    wire [7:0]  memDataRead, romRead, ramRead;
    wire [7:0]  memDataWrite;
    wire        memWrite;
    wire        memStrobe, romStrobe, ramStrobe;
    wire        romEnable, ramEnable;

    // 8k
    Memory #(.addrBusWidth(13)) rom(
        .clk(clk),
        .addr(memAddr[12:0]),
        .dataOut(romRead),
        .dataIn(memDataWrite),
        .write(1'b0),
        .strobe(romStrobe)
    );

    // 2k
    Memory #(.addrBusWidth(11)) ram(
        .clk(clk),
        .addr(memAddr[10:0]),
        .dataOut(ramRead),
        .dataIn(memDataWrite),
        .write(memWrite),
        .strobe(ramStrobe)
    );

    assign romEnable = memAddr[15] == 1'b0;
    assign ramEnable = memAddr[15] == 1'b1;
    assign romStrobe = memStrobe  & romEnable;
    assign ramStrobe = memStrobe  & ramEnable;
    assign memDataRead = romEnable ? romRead : ramRead;

    Processor proc(
        .clk(clk),
        .memAddr(memAddr),
        .memDataRead(memDataRead),
        .memDataWrite(memDataWrite),
        .memWrite(memWrite),
        .memStrobe(memStrobe),
        .port2Out(port2),
        .port3Out(port3)
    );
endmodule
