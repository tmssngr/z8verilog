localparam P01M = 8'hF8;
localparam FLAGS = 8'hFC;
localparam RP = 8'hFD;
localparam SPH = 8'hFE;
localparam SPL = 8'hFF;