localparam FLAG_INDEX_C = 7;
localparam FLAG_INDEX_Z = 6;
localparam FLAG_INDEX_S = 5;
localparam FLAG_INDEX_V = 4;
localparam FLAG_INDEX_D = 3; // 1 after sub, 0 after add
localparam FLAG_INDEX_H = 2; // half-carry

localparam FLAG_NONE = 0;
localparam FLAG_C = 8'h80;
localparam FLAG_Z = 8'h40;
localparam FLAG_S = 8'h20;
localparam FLAG_V = 8'h10;
localparam FLAG_D = 8'h08;
localparam FLAG_H = 8'h04;
