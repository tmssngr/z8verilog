localparam SIO   = 8'hF0;
localparam TMR   = 8'hF1;
localparam T1    = 8'hF2;
localparam PRE1  = 8'hF3;
localparam T0    = 8'hF4;
localparam PRE0  = 8'hF5;
localparam P3M   = 8'hF7;
localparam P01M  = 8'hF8;
localparam IPR   = 8'hF9;
localparam IRQ   = 8'hFA;
localparam IMR   = 8'hFB;
localparam FLAGS = 8'hFC;
localparam RP    = 8'hFD;
localparam SPH   = 8'hFE;
localparam SPL   = 8'hFF;
