localparam FETCH_MSB = 3;
localparam FETCH_INC  = 4'b1;
localparam FETCH_INSTR_WAIT  = 0;
localparam FETCH_INSTR_READ  = FETCH_INSTR_WAIT + 1;
localparam FETCH_SECOND_WAIT = FETCH_INSTR_READ + 1;
localparam FETCH_SECOND_READ = FETCH_SECOND_WAIT + 1;
localparam FETCH_THIRD_WAIT  = FETCH_SECOND_READ + 1;
localparam FETCH_THIRD_READ  = FETCH_THIRD_WAIT + 1;
localparam FETCH_DECODE      = FETCH_THIRD_READ + 1;

localparam OP_MSB = 3;
localparam OP_UNDECIDED = 0;
localparam OP_LD        = OP_UNDECIDED + 1;
localparam OP_ALU1      = OP_LD + 1;
localparam OP_ALU1WORD  = OP_ALU1 + 1;
localparam OP_ALU2      = OP_ALU1WORD + 1;
localparam OP_POP       = OP_ALU2 + 1;
localparam OP_PUSH_I    = OP_POP + 1;
localparam OP_PUSH_E    = OP_PUSH_I + 1;
localparam OP_DJNZ      = OP_PUSH_E + 1;
localparam OP_JP        = OP_DJNZ + 1;
localparam OP_CALL      = OP_JP + 1;
localparam OP_RET       = OP_CALL + 1;
localparam OP_IRET      = OP_RET + 1;
localparam OP_LDC       = OP_IRET + 1;
localparam OP_ILLEGAL   = OP_LDC + 1;

localparam OPSTATE_MSB = 2;
localparam OPSTATE_INC = 3'b1;
localparam OPSTATE0 = 0;
localparam OPSTATE1 = OPSTATE0 + 1;
localparam OPSTATE2 = OPSTATE1 + 1;
localparam OPSTATE3 = OPSTATE2 + 1;
localparam OPSTATE4 = OPSTATE3 + 1;
localparam OPSTATE5 = OPSTATE4 + 1;
localparam OPSTATE6 = OPSTATE5 + 1;
