memory[16'h0000] = 8'h08;
memory[16'h0001] = 8'h00;
memory[16'h0002] = 8'h08;
memory[16'h0003] = 8'h03;
memory[16'h0004] = 8'h08;
memory[16'h0005] = 8'h06;
memory[16'h0006] = 8'h08;
memory[16'h0007] = 8'h09;
memory[16'h0008] = 8'h08;
memory[16'h0009] = 8'h0c;
memory[16'h000a] = 8'h08;
memory[16'h000b] = 8'h0f;
memory[16'h000c] = 8'h31;
memory[16'h000d] = 8'h00;
memory[16'h000e] = 8'h3c;
memory[16'h000f] = 8'h0f;
memory[16'h0010] = 8'hff;
memory[16'h0011] = 8'h76;
memory[16'h0012] = 8'he3;
memory[16'h0013] = 8'h04;
memory[16'h0014] = 8'h3c;
memory[16'h0015] = 8'hff;
memory[16'h0016] = 8'heb;
memory[16'h0017] = 8'h05;
memory[16'h0018] = 8'h76;
memory[16'h0019] = 8'he3;
memory[16'h001a] = 8'h04;
memory[16'h001b] = 8'heb;
memory[16'h001c] = 8'h20;
memory[16'h001d] = 8'he6;
memory[16'h001e] = 8'hf8;
memory[16'h001f] = 8'hb6;
memory[16'h0020] = 8'he6;
memory[16'h0021] = 8'hf7;
memory[16'h0022] = 8'h08;
memory[16'h0023] = 8'h4c;
memory[16'h0024] = 8'h08;
memory[16'h0025] = 8'h5c;
memory[16'h0026] = 8'h12;
memory[16'h0027] = 8'hc2;
memory[16'h0028] = 8'h64;
memory[16'h0029] = 8'h60;
memory[16'h002a] = 8'he6;
memory[16'h002b] = 8'hd2;
memory[16'h002c] = 8'h64;
memory[16'h002d] = 8'hc2;
memory[16'h002e] = 8'h74;
memory[16'h002f] = 8'h60;
memory[16'h0030] = 8'he6;
memory[16'h0031] = 8'hd2;
memory[16'h0032] = 8'h64;
memory[16'h0033] = 8'hb2;
memory[16'h0034] = 8'h67;
memory[16'h0035] = 8'h31;
memory[16'h0036] = 8'hf0;
memory[16'h0037] = 8'hed;
memory[16'h0038] = 8'he0;
memory[16'h0039] = 8'h00;
memory[16'h003a] = 8'h8d;
memory[16'h003b] = 8'h08;
memory[16'h003c] = 8'h12;
memory[16'h003d] = 8'he6;
memory[16'h003e] = 8'hf8;
memory[16'h003f] = 8'h04;
memory[16'h0040] = 8'he6;
memory[16'h0041] = 8'hf1;
memory[16'h0042] = 8'hc0;
memory[16'h0043] = 8'h0c;
memory[16'h0044] = 8'hff;
memory[16'h0045] = 8'h1c;
memory[16'h0046] = 8'hff;
memory[16'h0047] = 8'hcf;
memory[16'h0048] = 8'h56;
memory[16'h0049] = 8'he3;
memory[16'h004a] = 8'hdf;
memory[16'h004b] = 8'h46;
memory[16'h004c] = 8'he3;
memory[16'h004d] = 8'h20;
memory[16'h004e] = 8'h10;
memory[16'h004f] = 8'he1;
memory[16'h0050] = 8'h10;
memory[16'h0051] = 8'he0;
memory[16'h0052] = 8'h76;
memory[16'h0053] = 8'he3;
memory[16'h0054] = 8'h04;
memory[16'h0055] = 8'h6b;
memory[16'h0056] = 8'h04;
memory[16'h0057] = 8'h7b;
memory[16'h0058] = 8'hf5;
memory[16'h0059] = 8'h8b;
memory[16'h005a] = 8'hed;
memory[16'h005b] = 8'he6;
memory[16'h005c] = 8'hf8;
memory[16'h005d] = 8'h7f;
memory[16'h005e] = 8'h8b;
memory[16'h005f] = 8'hfe;
memory[16'h0060] = 8'h46;
memory[16'h0061] = 8'h7f;
memory[16'h0062] = 8'h18;
memory[16'h0063] = 8'he4;
memory[16'h0064] = 8'h7f;
memory[16'h0065] = 8'hf8;
memory[16'h0066] = 8'h56;
memory[16'h0067] = 8'h03;
memory[16'h0068] = 8'hdf;
memory[16'h0069] = 8'h76;
memory[16'h006a] = 8'h03;
memory[16'h006b] = 8'h04;
memory[16'h006c] = 8'h6b;
memory[16'h006d] = 8'hfb;
memory[16'h006e] = 8'h56;
memory[16'h006f] = 8'h7f;
memory[16'h0070] = 8'hf7;
memory[16'h0071] = 8'h46;
memory[16'h0072] = 8'h03;
memory[16'h0073] = 8'h20;
memory[16'h0074] = 8'he4;
memory[16'h0075] = 8'h7f;
memory[16'h0076] = 8'hf8;
memory[16'h0077] = 8'hff;
memory[16'h0078] = 8'hbf;
memory[16'h0079] = 8'h28;
memory[16'h007a] = 8'he4;
memory[16'h007b] = 8'h38;
memory[16'h007c] = 8'he5;
memory[16'h007d] = 8'haf;
memory[16'h007e] = 8'h02;
memory[16'h007f] = 8'h35;
memory[16'h0080] = 8'h12;
memory[16'h0081] = 8'h24;
memory[16'h0082] = 8'h4b;
memory[16'h0083] = 8'h16;
memory[16'h0084] = 8'haf;
memory[16'h0085] = 8'h22;
memory[16'h0086] = 8'h35;
memory[16'h0087] = 8'h32;
memory[16'h0088] = 8'h24;
memory[16'h0089] = 8'h4b;
memory[16'h008a] = 8'h0f;
memory[16'h008b] = 8'haf;
memory[16'h008c] = 8'h76;
memory[16'h008d] = 8'he4;
memory[16'h008e] = 8'h80;
memory[16'h008f] = 8'h6b;
memory[16'h0090] = 8'he8;
memory[16'h0091] = 8'hb0;
memory[16'h0092] = 8'he2;
memory[16'h0093] = 8'hb0;
memory[16'h0094] = 8'he3;
memory[16'h0095] = 8'h8b;
memory[16'h0096] = 8'hee;
memory[16'h0097] = 8'h46;
memory[16'h0098] = 8'h0f;
memory[16'h0099] = 8'h80;
memory[16'h009a] = 8'h46;
memory[16'h009b] = 8'h0e;
memory[16'h009c] = 8'h80;
memory[16'h009d] = 8'haf;
memory[16'h009e] = 8'h88;
memory[16'h009f] = 8'he2;
memory[16'h00a0] = 8'hb2;
memory[16'h00a1] = 8'h84;
memory[16'h00a2] = 8'h9c;
memory[16'h00a3] = 8'h02;
memory[16'h00a4] = 8'h68;
memory[16'h00a5] = 8'he2;
memory[16'h00a6] = 8'h78;
memory[16'h00a7] = 8'he3;
memory[16'h00a8] = 8'hd6;
memory[16'h00a9] = 8'h00;
memory[16'h00aa] = 8'h8c;
memory[16'h00ab] = 8'h48;
memory[16'h00ac] = 8'he6;
memory[16'h00ad] = 8'h58;
memory[16'h00ae] = 8'he7;
memory[16'h00af] = 8'h9a;
memory[16'h00b0] = 8'hf3;
memory[16'h00b1] = 8'h68;
memory[16'h00b2] = 8'he2;
memory[16'h00b3] = 8'h78;
memory[16'h00b4] = 8'he3;
memory[16'h00b5] = 8'hb0;
memory[16'h00b6] = 8'he2;
memory[16'h00b7] = 8'hb0;
memory[16'h00b8] = 8'he3;
memory[16'h00b9] = 8'haf;
memory[16'h00ba] = 8'hd6;
memory[16'h00bb] = 8'h00;
memory[16'h00bc] = 8'h9e;
memory[16'h00bd] = 8'hbc;
memory[16'h00be] = 8'h0f;
memory[16'h00bf] = 8'hd0;
memory[16'h00c0] = 8'he6;
memory[16'h00c1] = 8'hc0;
memory[16'h00c2] = 8'he7;
memory[16'h00c3] = 8'hfb;
memory[16'h00c4] = 8'h06;
memory[16'h00c5] = 8'h02;
memory[16'h00c6] = 8'h35;
memory[16'h00c7] = 8'h12;
memory[16'h00c8] = 8'h24;
memory[16'h00c9] = 8'h4b;
memory[16'h00ca] = 8'hcc;
memory[16'h00cb] = 8'h10;
memory[16'h00cc] = 8'he5;
memory[16'h00cd] = 8'h10;
memory[16'h00ce] = 8'he4;
memory[16'h00cf] = 8'hcb;
memory[16'h00d0] = 8'h04;
memory[16'h00d1] = 8'h42;
memory[16'h00d2] = 8'h67;
memory[16'h00d3] = 8'heb;
memory[16'h00d4] = 8'hc2;
memory[16'h00d5] = 8'hba;
memory[16'h00d6] = 8'he8;
memory[16'h00d7] = 8'h48;
memory[16'h00d8] = 8'he2;
memory[16'h00d9] = 8'h58;
memory[16'h00da] = 8'he3;
memory[16'h00db] = 8'h10;
memory[16'h00dc] = 8'he8;
memory[16'h00dd] = 8'h7b;
memory[16'h00de] = 8'hb2;
memory[16'h00df] = 8'haf;
memory[16'h00e0] = 8'hd6;
memory[16'h00e1] = 8'h00;
memory[16'h00e2] = 8'h9e;
memory[16'h00e3] = 8'h9c;
memory[16'h00e4] = 8'h10;
memory[16'h00e5] = 8'hcf;
memory[16'h00e6] = 8'hb0;
memory[16'h00e7] = 8'hea;
memory[16'h00e8] = 8'hb0;
memory[16'h00e9] = 8'heb;
memory[16'h00ea] = 8'h10;
memory[16'h00eb] = 8'he7;
memory[16'h00ec] = 8'h10;
memory[16'h00ed] = 8'he6;
memory[16'h00ee] = 8'h10;
memory[16'h00ef] = 8'heb;
memory[16'h00f0] = 8'h10;
memory[16'h00f1] = 8'hea;
memory[16'h00f2] = 8'h7b;
memory[16'h00f3] = 8'h0a;
memory[16'h00f4] = 8'ha2;
memory[16'h00f5] = 8'h4a;
memory[16'h00f6] = 8'hbb;
memory[16'h00f7] = 8'h0b;
memory[16'h00f8] = 8'h7b;
memory[16'h00f9] = 8'h04;
memory[16'h00fa] = 8'ha2;
memory[16'h00fb] = 8'h5b;
memory[16'h00fc] = 8'hbb;
memory[16'h00fd] = 8'h05;
memory[16'h00fe] = 8'h22;
memory[16'h00ff] = 8'hb5;
memory[16'h0100] = 8'h32;
memory[16'h0101] = 8'ha4;
memory[16'h0102] = 8'hdf;
memory[16'h0103] = 8'h9a;
memory[16'h0104] = 8'he5;
memory[16'h0105] = 8'h98;
memory[16'h0106] = 8'he4;
memory[16'h0107] = 8'h42;
memory[16'h0108] = 8'h95;
memory[16'h0109] = 8'h6b;
memory[16'h010a] = 8'h0a;
memory[16'h010b] = 8'h10;
memory[16'h010c] = 8'he7;
memory[16'h010d] = 8'h10;
memory[16'h010e] = 8'he6;
memory[16'h010f] = 8'h28;
memory[16'h0110] = 8'he6;
memory[16'h0111] = 8'h38;
memory[16'h0112] = 8'he7;
memory[16'h0113] = 8'h8b;
memory[16'h0114] = 8'hc2;
memory[16'h0115] = 8'hd6;
memory[16'h0116] = 8'h01;
memory[16'h0117] = 8'h0f;
memory[16'h0118] = 8'h46;
memory[16'h0119] = 8'h0e;
memory[16'h011a] = 8'h40;
memory[16'h011b] = 8'h46;
memory[16'h011c] = 8'h0f;
memory[16'h011d] = 8'h80;
memory[16'h011e] = 8'haf;
memory[16'h011f] = 8'hd6;
memory[16'h0120] = 8'h00;
memory[16'h0121] = 8'he0;
memory[16'h0122] = 8'h88;
memory[16'h0123] = 8'he2;
memory[16'h0124] = 8'h28;
memory[16'h0125] = 8'hea;
memory[16'h0126] = 8'h38;
memory[16'h0127] = 8'heb;
memory[16'h0128] = 8'h8b;
memory[16'h0129] = 8'had;
memory[16'h012a] = 8'h42;
memory[16'h012b] = 8'h24;
memory[16'h012c] = 8'h42;
memory[16'h012d] = 8'h35;
memory[16'h012e] = 8'haf;
memory[16'h012f] = 8'h52;
memory[16'h0130] = 8'h24;
memory[16'h0131] = 8'h52;
memory[16'h0132] = 8'h35;
memory[16'h0133] = 8'haf;
memory[16'h0134] = 8'hb2;
memory[16'h0135] = 8'h24;
memory[16'h0136] = 8'hb2;
memory[16'h0137] = 8'h35;
memory[16'h0138] = 8'haf;
memory[16'h0139] = 8'hd6;
memory[16'h013a] = 8'h00;
memory[16'h013b] = 8'h79;
memory[16'h013c] = 8'h60;
memory[16'h013d] = 8'he2;
memory[16'h013e] = 8'h60;
memory[16'h013f] = 8'he3;
memory[16'h0140] = 8'haf;
memory[16'h0141] = 8'h56;
memory[16'h0142] = 8'h0f;
memory[16'h0143] = 8'h8f;
memory[16'h0144] = 8'ha2;
memory[16'h0145] = 8'h24;
memory[16'h0146] = 8'h6b;
memory[16'h0147] = 8'h0a;
memory[16'h0148] = 8'h7c;
memory[16'h0149] = 8'h20;
memory[16'h014a] = 8'hab;
memory[16'h014b] = 8'h02;
memory[16'h014c] = 8'h7c;
memory[16'h014d] = 8'h10;
memory[16'h014e] = 8'h44;
memory[16'h014f] = 8'he7;
memory[16'h0150] = 8'h0f;
memory[16'h0151] = 8'haf;
memory[16'h0152] = 8'h7c;
memory[16'h0153] = 8'h40;
memory[16'h0154] = 8'ha2;
memory[16'h0155] = 8'h35;
memory[16'h0156] = 8'h6b;
memory[16'h0157] = 8'hf6;
memory[16'h0158] = 8'h7c;
memory[16'h0159] = 8'h20;
memory[16'h015a] = 8'hbb;
memory[16'h015b] = 8'hf2;
memory[16'h015c] = 8'h8b;
memory[16'h015d] = 8'hee;
memory[16'h015e] = 8'h88;
memory[16'h015f] = 8'he3;
memory[16'h0160] = 8'h78;
memory[16'h0161] = 8'he3;
memory[16'h0162] = 8'h68;
memory[16'h0163] = 8'he2;
memory[16'h0164] = 8'h58;
memory[16'h0165] = 8'he2;
memory[16'h0166] = 8'hf0;
memory[16'h0167] = 8'he5;
memory[16'h0168] = 8'hf0;
memory[16'h0169] = 8'he7;
memory[16'h016a] = 8'h4c;
memory[16'h016b] = 8'h25;
memory[16'h016c] = 8'hac;
memory[16'h016d] = 8'h04;
memory[16'h016e] = 8'hbc;
memory[16'h016f] = 8'h15;
memory[16'h0170] = 8'h57;
memory[16'h0171] = 8'heb;
memory[16'h0172] = 8'h0f;
memory[16'h0173] = 8'h07;
memory[16'h0174] = 8'heb;
memory[16'h0175] = 8'h30;
memory[16'h0176] = 8'ha7;
memory[16'h0177] = 8'heb;
memory[16'h0178] = 8'h3a;
memory[16'h0179] = 8'h7b;
memory[16'h017a] = 8'h03;
memory[16'h017b] = 8'h07;
memory[16'h017c] = 8'heb;
memory[16'h017d] = 8'h07;
memory[16'h017e] = 8'hbe;
memory[16'h017f] = 8'haa;
memory[16'h0180] = 8'hef;
memory[16'h0181] = 8'haf;
memory[16'h0182] = 8'h48;
memory[16'h0183] = 8'he2;
memory[16'h0184] = 8'h58;
memory[16'h0185] = 8'he3;
memory[16'h0186] = 8'hd6;
memory[16'h0187] = 8'h00;
memory[16'h0188] = 8'h8c;
memory[16'h0189] = 8'h10;
memory[16'h018a] = 8'he4;
memory[16'h018b] = 8'h4c;
memory[16'h018c] = 8'h20;
memory[16'h018d] = 8'hfb;
memory[16'h018e] = 8'h02;
memory[16'h018f] = 8'h4c;
memory[16'h0190] = 8'h2d;
memory[16'h0191] = 8'hbc;
memory[16'h0192] = 8'h06;
memory[16'h0193] = 8'hac;
memory[16'h0194] = 8'h15;
memory[16'h0195] = 8'hb1;
memory[16'h0196] = 8'hea;
memory[16'h0197] = 8'hae;
memory[16'h0198] = 8'hba;
memory[16'h0199] = 8'hfb;
memory[16'h019a] = 8'hbc;
memory[16'h019b] = 8'h0f;
memory[16'h019c] = 8'hd0;
memory[16'h019d] = 8'he2;
memory[16'h019e] = 8'hc0;
memory[16'h019f] = 8'he3;
memory[16'h01a0] = 8'hfb;
memory[16'h01a1] = 8'h0c;
memory[16'h01a2] = 8'h02;
memory[16'h01a3] = 8'h7a;
memory[16'h01a4] = 8'h40;
memory[16'h01a5] = 8'he7;
memory[16'h01a6] = 8'h12;
memory[16'h01a7] = 8'h69;
memory[16'h01a8] = 8'h40;
memory[16'h01a9] = 8'he6;
memory[16'h01aa] = 8'h12;
memory[16'h01ab] = 8'h58;
memory[16'h01ac] = 8'h40;
memory[16'h01ad] = 8'he5;
memory[16'h01ae] = 8'h02;
memory[16'h01af] = 8'haa;
memory[16'h01b0] = 8'h40;
memory[16'h01b1] = 8'hea;
memory[16'h01b2] = 8'h12;
memory[16'h01b3] = 8'h99;
memory[16'h01b4] = 8'h40;
memory[16'h01b5] = 8'he9;
memory[16'h01b6] = 8'h12;
memory[16'h01b7] = 8'h88;
memory[16'h01b8] = 8'h40;
memory[16'h01b9] = 8'he8;
memory[16'h01ba] = 8'hba;
memory[16'h01bb] = 8'he0;
memory[16'h01bc] = 8'h88;
memory[16'h01bd] = 8'he7;
memory[16'h01be] = 8'h98;
memory[16'h01bf] = 8'he7;
memory[16'h01c0] = 8'h78;
memory[16'h01c1] = 8'he6;
memory[16'h01c2] = 8'hf0;
memory[16'h01c3] = 8'he6;
memory[16'h01c4] = 8'hf0;
memory[16'h01c5] = 8'he8;
memory[16'h01c6] = 8'hac;
memory[16'h01c7] = 8'h05;
memory[16'h01c8] = 8'h8b;
memory[16'h01c9] = 8'ha4;
memory[16'h01ca] = 8'hf1;
memory[16'h01cb] = 8'hed;
memory[16'h01cc] = 8'hec;
memory[16'h01cd] = 8'h04;
memory[16'h01ce] = 8'h11;
memory[16'h01cf] = 8'hed;
memory[16'h01d0] = 8'h10;
memory[16'h01d1] = 8'he5;
memory[16'h01d2] = 8'h10;
memory[16'h01d3] = 8'he4;
memory[16'h01d4] = 8'h10;
memory[16'h01d5] = 8'he3;
memory[16'h01d6] = 8'hea;
memory[16'h01d7] = 8'hf6;
memory[16'h01d8] = 8'haf;
memory[16'h01d9] = 8'hdc;
memory[16'h01da] = 8'h16;
memory[16'h01db] = 8'hb0;
memory[16'h01dc] = 8'he4;
memory[16'h01dd] = 8'hb0;
memory[16'h01de] = 8'he5;
memory[16'h01df] = 8'ha6;
memory[16'h01e0] = 8'he6;
memory[16'h01e1] = 8'h25;
memory[16'h01e2] = 8'heb;
memory[16'h01e3] = 8'h27;
memory[16'h01e4] = 8'hcc;
memory[16'h01e5] = 8'h05;
memory[16'h01e6] = 8'hde;
memory[16'h01e7] = 8'h27;
memory[16'h01e8] = 8'hed;
memory[16'h01e9] = 8'h30;
memory[16'h01ea] = 8'h7b;
memory[16'h01eb] = 8'h19;
memory[16'h01ec] = 8'ha7;
memory[16'h01ed] = 8'hed;
memory[16'h01ee] = 8'h0a;
memory[16'h01ef] = 8'h7b;
memory[16'h01f0] = 8'h0d;
memory[16'h01f1] = 8'h27;
memory[16'h01f2] = 8'hed;
memory[16'h01f3] = 8'h11;
memory[16'h01f4] = 8'h7b;
memory[16'h01f5] = 8'h0f;
memory[16'h01f6] = 8'h07;
memory[16'h01f7] = 8'hed;
memory[16'h01f8] = 8'h0a;
memory[16'h01f9] = 8'ha7;
memory[16'h01fa] = 8'hed;
memory[16'h01fb] = 8'h10;
memory[16'h01fc] = 8'hfb;
memory[16'h01fd] = 8'h07;
memory[16'h01fe] = 8'hd6;
memory[16'h01ff] = 8'h01;
memory[16'h0200] = 8'hca;
memory[16'h0201] = 8'hca;
memory[16'h0202] = 8'he3;
memory[16'h0203] = 8'hcf;
memory[16'h0204] = 8'haf;
memory[16'h0205] = 8'ha6;
memory[16'h0206] = 8'hec;
memory[16'h0207] = 8'h05;
memory[16'h0208] = 8'h6b;
memory[16'h0209] = 8'hf9;
memory[16'h020a] = 8'haf;
memory[16'h020b] = 8'hcc;
memory[16'h020c] = 8'h06;
memory[16'h020d] = 8'hb0;
memory[16'h020e] = 8'he2;
memory[16'h020f] = 8'hb0;
memory[16'h0210] = 8'he3;
memory[16'h0211] = 8'ha6;
memory[16'h0212] = 8'he6;
memory[16'h0213] = 8'h2d;
memory[16'h0214] = 8'heb;
memory[16'h0215] = 8'h02;
memory[16'h0216] = 8'h2e;
memory[16'h0217] = 8'hde;
memory[16'h0218] = 8'h27;
memory[16'h0219] = 8'hed;
memory[16'h021a] = 8'h30;
memory[16'h021b] = 8'h7b;
memory[16'h021c] = 8'h0c;
memory[16'h021d] = 8'ha7;
memory[16'h021e] = 8'hed;
memory[16'h021f] = 8'h0a;
memory[16'h0220] = 8'hfb;
memory[16'h0221] = 8'h07;
memory[16'h0222] = 8'hd6;
memory[16'h0223] = 8'h01;
memory[16'h0224] = 8'hca;
memory[16'h0225] = 8'hca;
memory[16'h0226] = 8'hf0;
memory[16'h0227] = 8'hcf;
memory[16'h0228] = 8'haf;
memory[16'h0229] = 8'ha6;
memory[16'h022a] = 8'hec;
memory[16'h022b] = 8'h06;
memory[16'h022c] = 8'h6b;
memory[16'h022d] = 8'hf9;
memory[16'h022e] = 8'ha6;
memory[16'h022f] = 8'he3;
memory[16'h0230] = 8'h04;
memory[16'h0231] = 8'hfb;
memory[16'h0232] = 8'hf4;
memory[16'h0233] = 8'hb0;
memory[16'h0234] = 8'he6;
memory[16'h0235] = 8'hb0;
memory[16'h0236] = 8'he7;
memory[16'h0237] = 8'hbc;
memory[16'h0238] = 8'h13;
memory[16'h0239] = 8'h8c;
memory[16'h023a] = 8'h27;
memory[16'h023b] = 8'h9c;
memory[16'h023c] = 8'h10;
memory[16'h023d] = 8'hd6;
memory[16'h023e] = 8'h02;
memory[16'h023f] = 8'h71;
memory[16'h0240] = 8'hbe;
memory[16'h0241] = 8'h8c;
memory[16'h0242] = 8'h03;
memory[16'h0243] = 8'h9c;
memory[16'h0244] = 8'he8;
memory[16'h0245] = 8'hd6;
memory[16'h0246] = 8'h02;
memory[16'h0247] = 8'h6f;
memory[16'h0248] = 8'h8c;
memory[16'h0249] = 8'h00;
memory[16'h024a] = 8'h9c;
memory[16'h024b] = 8'h64;
memory[16'h024c] = 8'hd6;
memory[16'h024d] = 8'h02;
memory[16'h024e] = 8'h6f;
memory[16'h024f] = 8'hbe;
memory[16'h0250] = 8'h9c;
memory[16'h0251] = 8'h0a;
memory[16'h0252] = 8'hd6;
memory[16'h0253] = 8'h02;
memory[16'h0254] = 8'h6f;
memory[16'h0255] = 8'h9c;
memory[16'h0256] = 8'h01;
memory[16'h0257] = 8'hd6;
memory[16'h0258] = 8'h02;
memory[16'h0259] = 8'h6f;
memory[16'h025a] = 8'h48;
memory[16'h025b] = 8'he6;
memory[16'h025c] = 8'h58;
memory[16'h025d] = 8'he7;
memory[16'h025e] = 8'h10;
memory[16'h025f] = 8'he6;
memory[16'h0260] = 8'h7b;
memory[16'h0261] = 8'hc5;
memory[16'h0262] = 8'hc0;
memory[16'h0263] = 8'he2;
memory[16'h0264] = 8'hfb;
memory[16'h0265] = 8'h18;
memory[16'h0266] = 8'hd6;
memory[16'h0267] = 8'h00;
memory[16'h0268] = 8'h91;
memory[16'h0269] = 8'h48;
memory[16'h026a] = 8'he2;
memory[16'h026b] = 8'h58;
memory[16'h026c] = 8'he3;
memory[16'h026d] = 8'h8b;
memory[16'h026e] = 8'h0f;
memory[16'h026f] = 8'hf1;
memory[16'h0270] = 8'heb;
memory[16'h0271] = 8'he3;
memory[16'h0272] = 8'hab;
memory[16'h0273] = 8'h56;
memory[16'h0274] = 8'hea;
memory[16'h0275] = 8'h0f;
memory[16'h0276] = 8'h6b;
memory[16'h0277] = 8'h06;
memory[16'h0278] = 8'h02;
memory[16'h0279] = 8'h79;
memory[16'h027a] = 8'h12;
memory[16'h027b] = 8'h68;
memory[16'h027c] = 8'haa;
memory[16'h027d] = 8'hfa;
memory[16'h027e] = 8'hdf;
memory[16'h027f] = 8'haf;
memory[16'h0280] = 8'h50;
memory[16'h0281] = 8'he8;
memory[16'h0282] = 8'h50;
memory[16'h0283] = 8'he9;
memory[16'h0284] = 8'h50;
memory[16'h0285] = 8'he2;
memory[16'h0286] = 8'h50;
memory[16'h0287] = 8'he3;
memory[16'h0288] = 8'h50;
memory[16'h0289] = 8'he6;
memory[16'h028a] = 8'h50;
memory[16'h028b] = 8'he7;
memory[16'h028c] = 8'h30;
memory[16'h028d] = 8'he8;
memory[16'h028e] = 8'hd6;
memory[16'h028f] = 8'h02;
memory[16'h0290] = 8'h80;
memory[16'h0291] = 8'hf3;
memory[16'h0292] = 8'h74;
memory[16'h0293] = 8'h7e;
memory[16'h0294] = 8'h8b;
memory[16'h0295] = 8'h03;
memory[16'h0296] = 8'hd6;
memory[16'h0297] = 8'h02;
memory[16'h0298] = 8'h80;
memory[16'h0299] = 8'hf3;
memory[16'h029a] = 8'h75;
memory[16'h029b] = 8'h30;
memory[16'h029c] = 8'he2;
memory[16'h029d] = 8'hd6;
memory[16'h029e] = 8'h02;
memory[16'h029f] = 8'h80;
memory[16'h02a0] = 8'h92;
memory[16'h02a1] = 8'h46;
memory[16'h02a2] = 8'ha0;
memory[16'h02a3] = 8'he6;
memory[16'h02a4] = 8'h8b;
memory[16'h02a5] = 8'h03;
memory[16'h02a6] = 8'hd6;
memory[16'h02a7] = 8'h02;
memory[16'h02a8] = 8'h80;
memory[16'h02a9] = 8'h92;
memory[16'h02aa] = 8'h56;
memory[16'h02ab] = 8'h30;
memory[16'h02ac] = 8'he2;
memory[16'h02ad] = 8'he3;
memory[16'h02ae] = 8'h25;
memory[16'h02af] = 8'h5e;
memory[16'h02b0] = 8'h0d;
memory[16'h02b1] = 8'hb0;
memory[16'h02b2] = 8'he2;
memory[16'h02b3] = 8'he3;
memory[16'h02b4] = 8'h35;
memory[16'h02b5] = 8'haf;
memory[16'h02b6] = 8'h82;
memory[16'h02b7] = 8'h24;
memory[16'h02b8] = 8'ha0;
memory[16'h02b9] = 8'he4;
memory[16'h02ba] = 8'h0d;
memory[16'h02bb] = 8'hb0;
memory[16'h02bc] = 8'he2;
memory[16'h02bd] = 8'h82;
memory[16'h02be] = 8'h34;
memory[16'h02bf] = 8'haf;
memory[16'h02c0] = 8'hd6;
memory[16'h02c1] = 8'h02;
memory[16'h02c2] = 8'hc8;
memory[16'h02c3] = 8'h5c;
memory[16'h02c4] = 8'h20;
memory[16'h02c5] = 8'hd6;
memory[16'h02c6] = 8'h08;
memory[16'h02c7] = 8'h18;
memory[16'h02c8] = 8'h5c;
memory[16'h02c9] = 8'h08;
memory[16'h02ca] = 8'h8d;
memory[16'h02cb] = 8'h08;
memory[16'h02cc] = 8'h18;
memory[16'h02cd] = 8'hcf;
memory[16'h02ce] = 8'h10;
memory[16'h02cf] = 8'he5;
memory[16'h02d0] = 8'h10;
memory[16'h02d1] = 8'he4;
memory[16'h02d2] = 8'h16;
memory[16'h02d3] = 8'he5;
memory[16'h02d4] = 8'h00;
memory[16'h02d5] = 8'h8d;
memory[16'h02d6] = 8'h00;
memory[16'h02d7] = 8'h79;
memory[16'h02d8] = 8'hcf;
memory[16'h02d9] = 8'hc0;
memory[16'h02da] = 8'he4;
memory[16'h02db] = 8'hc0;
memory[16'h02dc] = 8'he5;
memory[16'h02dd] = 8'hfb;
memory[16'h02de] = 8'hf6;
memory[16'h02df] = 8'h46;
memory[16'h02e0] = 8'he4;
memory[16'h02e1] = 8'h80;
memory[16'h02e2] = 8'h8b;
memory[16'h02e3] = 8'hf1;
memory[16'h02e4] = 8'h5c;
memory[16'h02e5] = 8'h3f;
memory[16'h02e6] = 8'hd6;
memory[16'h02e7] = 8'h08;
memory[16'h02e8] = 8'h18;
memory[16'h02e9] = 8'hfc;
memory[16'h02ea] = 8'h15;
memory[16'h02eb] = 8'hfe;
memory[16'h02ec] = 8'ha6;
memory[16'h02ed] = 8'hef;
memory[16'h02ee] = 8'h1f;
memory[16'h02ef] = 8'h6b;
memory[16'h02f0] = 8'h20;
memory[16'h02f1] = 8'hd6;
memory[16'h02f2] = 8'h08;
memory[16'h02f3] = 8'h15;
memory[16'h02f4] = 8'hf3;
memory[16'h02f5] = 8'hf3;
memory[16'h02f6] = 8'ha6;
memory[16'h02f7] = 8'he3;
memory[16'h02f8] = 8'h0d;
memory[16'h02f9] = 8'h6b;
memory[16'h02fa] = 8'h16;
memory[16'h02fb] = 8'ha6;
memory[16'h02fc] = 8'he3;
memory[16'h02fd] = 8'h08;
memory[16'h02fe] = 8'heb;
memory[16'h02ff] = 8'h19;
memory[16'h0300] = 8'h5c;
memory[16'h0301] = 8'h20;
memory[16'h0302] = 8'hd6;
memory[16'h0303] = 8'h08;
memory[16'h0304] = 8'h18;
memory[16'h0305] = 8'h00;
memory[16'h0306] = 8'hef;
memory[16'h0307] = 8'ha6;
memory[16'h0308] = 8'hef;
memory[16'h0309] = 8'h15;
memory[16'h030a] = 8'h6b;
memory[16'h030b] = 8'hdf;
memory[16'h030c] = 8'hd6;
memory[16'h030d] = 8'h02;
memory[16'h030e] = 8'hc8;
memory[16'h030f] = 8'h8b;
memory[16'h0310] = 8'he0;
memory[16'h0311] = 8'hd6;
memory[16'h0312] = 8'h01;
memory[16'h0313] = 8'hd9;
memory[16'h0314] = 8'hfb;
memory[16'h0315] = 8'hce;
memory[16'h0316] = 8'h8d;
memory[16'h0317] = 8'h00;
memory[16'h0318] = 8'h79;
memory[16'h0319] = 8'h3e;
memory[16'h031a] = 8'hdb;
memory[16'h031b] = 8'hcf;
memory[16'h031c] = 8'ha6;
memory[16'h031d] = 8'hef;
memory[16'h031e] = 8'h16;
memory[16'h031f] = 8'h6b;
memory[16'h0320] = 8'hc8;
memory[16'h0321] = 8'hd6;
memory[16'h0322] = 8'h02;
memory[16'h0323] = 8'hc0;
memory[16'h0324] = 8'h00;
memory[16'h0325] = 8'hef;
memory[16'h0326] = 8'h8b;
memory[16'h0327] = 8'hf4;
memory[16'h0328] = 8'h03;
memory[16'h0329] = 8'h4e;
memory[16'h032a] = 8'h4f;
memory[16'h032b] = 8'h54;
memory[16'h032c] = 8'h01;
memory[16'h032d] = 8'h39;
memory[16'h032e] = 8'h03;
memory[16'h032f] = 8'h41;
memory[16'h0330] = 8'h42;
memory[16'h0331] = 8'h53;
memory[16'h0332] = 8'h00;
memory[16'h0333] = 8'h8c;
memory[16'h0334] = 8'h05;
memory[16'h0335] = 8'h53;
memory[16'h0336] = 8'h45;
memory[16'h0337] = 8'h54;
memory[16'h0338] = 8'h52;
memory[16'h0339] = 8'h52;
memory[16'h033a] = 8'h02;
memory[16'h033b] = 8'h8e;
memory[16'h033c] = 8'h04;
memory[16'h033d] = 8'h53;
memory[16'h033e] = 8'h45;
memory[16'h033f] = 8'h54;
memory[16'h0340] = 8'h52;
memory[16'h0341] = 8'h02;
memory[16'h0342] = 8'h96;
memory[16'h0343] = 8'h05;
memory[16'h0344] = 8'h53;
memory[16'h0345] = 8'h45;
memory[16'h0346] = 8'h54;
memory[16'h0347] = 8'h45;
memory[16'h0348] = 8'h57;
memory[16'h0349] = 8'h02;
memory[16'h034a] = 8'h9d;
memory[16'h034b] = 8'h05;
memory[16'h034c] = 8'h53;
memory[16'h034d] = 8'h45;
memory[16'h034e] = 8'h54;
memory[16'h034f] = 8'h45;
memory[16'h0350] = 8'h42;
memory[16'h0351] = 8'h02;
memory[16'h0352] = 8'ha6;
memory[16'h0353] = 8'h05;
memory[16'h0354] = 8'h47;
memory[16'h0355] = 8'h45;
memory[16'h0356] = 8'h54;
memory[16'h0357] = 8'h52;
memory[16'h0358] = 8'h52;
memory[16'h0359] = 8'h02;
memory[16'h035a] = 8'had;
memory[16'h035b] = 8'h04;
memory[16'h035c] = 8'h47;
memory[16'h035d] = 8'h45;
memory[16'h035e] = 8'h54;
memory[16'h035f] = 8'h52;
memory[16'h0360] = 8'h02;
memory[16'h0361] = 8'hb1;
memory[16'h0362] = 8'h05;
memory[16'h0363] = 8'h47;
memory[16'h0364] = 8'h45;
memory[16'h0365] = 8'h54;
memory[16'h0366] = 8'h45;
memory[16'h0367] = 8'h57;
memory[16'h0368] = 8'h02;
memory[16'h0369] = 8'hb6;
memory[16'h036a] = 8'h05;
memory[16'h036b] = 8'h47;
memory[16'h036c] = 8'h45;
memory[16'h036d] = 8'h54;
memory[16'h036e] = 8'h45;
memory[16'h036f] = 8'h42;
memory[16'h0370] = 8'h02;
memory[16'h0371] = 8'hbb;
memory[16'h0372] = 8'h02;
memory[16'h0373] = 8'h52;
memory[16'h0374] = 8'h4c;
memory[16'h0375] = 8'h02;
memory[16'h0376] = 8'hcd;
memory[16'h0377] = 8'h02;
memory[16'h0378] = 8'h52;
memory[16'h0379] = 8'h52;
memory[16'h037a] = 8'h02;
memory[16'h037b] = 8'hd8;
memory[16'h037c] = 8'h05;
memory[16'h037d] = 8'h49;
memory[16'h037e] = 8'h4e;
memory[16'h037f] = 8'h50;
memory[16'h0380] = 8'h55;
memory[16'h0381] = 8'h54;
memory[16'h0382] = 8'h02;
memory[16'h0383] = 8'he4;
memory[16'h0384] = 8'h03;
memory[16'h0385] = 8'h47;
memory[16'h0386] = 8'h54;
memory[16'h0387] = 8'h43;
memory[16'h0388] = 8'h08;
memory[16'h0389] = 8'h15;
memory[16'h038a] = 8'h03;
memory[16'h038b] = 8'h50;
memory[16'h038c] = 8'h54;
memory[16'h038d] = 8'h43;
memory[16'h038e] = 8'h08;
memory[16'h038f] = 8'h18;
memory[16'h0390] = 8'hff;
memory[16'h0391] = 8'hfc;
memory[16'h0392] = 8'h16;
memory[16'h0393] = 8'hc2;
memory[16'h0394] = 8'h60;
memory[16'h0395] = 8'ha0;
memory[16'h0396] = 8'he0;
memory[16'h0397] = 8'ha2;
memory[16'h0398] = 8'h67;
memory[16'h0399] = 8'haf;
memory[16'h039a] = 8'hac;
memory[16'h039b] = 8'h03;
memory[16'h039c] = 8'hbc;
memory[16'h039d] = 8'hc1;
memory[16'h039e] = 8'hdc;
memory[16'h039f] = 8'h03;
memory[16'h03a0] = 8'hd6;
memory[16'h03a1] = 8'h03;
memory[16'h03a2] = 8'haf;
memory[16'h03a3] = 8'h6b;
memory[16'h03a4] = 8'h1b;
memory[16'h03a5] = 8'ha6;
memory[16'h03a6] = 8'he6;
memory[16'h03a7] = 8'h24;
memory[16'h03a8] = 8'heb;
memory[16'h03a9] = 8'h16;
memory[16'h03aa] = 8'hd6;
memory[16'h03ab] = 8'h03;
memory[16'h03ac] = 8'h91;
memory[16'h03ad] = 8'hdc;
memory[16'h03ae] = 8'h03;
memory[16'h03af] = 8'hd6;
memory[16'h03b0] = 8'h03;
memory[16'h03b1] = 8'hb6;
memory[16'h03b2] = 8'h6b;
memory[16'h03b3] = 8'h0c;
memory[16'h03b4] = 8'hda;
memory[16'h03b5] = 8'hf9;
memory[16'h03b6] = 8'hcc;
memory[16'h03b7] = 8'h17;
memory[16'h03b8] = 8'hc3;
memory[16'h03b9] = 8'hca;
memory[16'h03ba] = 8'hc3;
memory[16'h03bb] = 8'hca;
memory[16'h03bc] = 8'hc3;
memory[16'h03bd] = 8'hca;
memory[16'h03be] = 8'ha2;
memory[16'h03bf] = 8'h67;
memory[16'h03c0] = 8'haf;
memory[16'h03c1] = 8'h2b;
memory[16'h03c2] = 8'h00;
memory[16'h03c3] = 8'h7e;
memory[16'h03c4] = 8'h2d;
memory[16'h03c5] = 8'h00;
memory[16'h03c6] = 8'h85;
memory[16'h03c7] = 8'h2a;
memory[16'h03c8] = 8'h00;
memory[16'h03c9] = 8'hba;
memory[16'h03ca] = 8'h2f;
memory[16'h03cb] = 8'h00;
memory[16'h03cc] = 8'he0;
memory[16'h03cd] = 8'h41;
memory[16'h03ce] = 8'h01;
memory[16'h03cf] = 8'h2f;
memory[16'h03d0] = 8'h4f;
memory[16'h03d1] = 8'h01;
memory[16'h03d2] = 8'h2a;
memory[16'h03d3] = 8'h58;
memory[16'h03d4] = 8'h01;
memory[16'h03d5] = 8'h34;
memory[16'h03d6] = 8'h4d;
memory[16'h03d7] = 8'h01;
memory[16'h03d8] = 8'h1f;
memory[16'h03d9] = 8'ha7;
memory[16'h03da] = 8'hef;
memory[16'h03db] = 8'h41;
memory[16'h03dc] = 8'h7b;
memory[16'h03dd] = 8'h12;
memory[16'h03de] = 8'ha7;
memory[16'h03df] = 8'hef;
memory[16'h03e0] = 8'h5b;
memory[16'h03e1] = 8'haf;
memory[16'h03e2] = 8'hd6;
memory[16'h03e3] = 8'h03;
memory[16'h03e4] = 8'hd9;
memory[16'h03e5] = 8'h7b;
memory[16'h03e6] = 8'h08;
memory[16'h03e7] = 8'ha7;
memory[16'h03e8] = 8'hef;
memory[16'h03e9] = 8'h30;
memory[16'h03ea] = 8'h7b;
memory[16'h03eb] = 8'h04;
memory[16'h03ec] = 8'ha7;
memory[16'h03ed] = 8'hef;
memory[16'h03ee] = 8'h3a;
memory[16'h03ef] = 8'haf;
memory[16'h03f0] = 8'hcf;
memory[16'h03f1] = 8'haf;
memory[16'h03f2] = 8'hd6;
memory[16'h03f3] = 8'h03;
memory[16'h03f4] = 8'he7;
memory[16'h03f5] = 8'h7b;
memory[16'h03f6] = 8'hf8;
memory[16'h03f7] = 8'ha7;
memory[16'h03f8] = 8'hef;
memory[16'h03f9] = 8'h41;
memory[16'h03fa] = 8'h7b;
memory[16'h03fb] = 8'hf4;
memory[16'h03fc] = 8'ha7;
memory[16'h03fd] = 8'hef;
memory[16'h03fe] = 8'h47;
memory[16'h03ff] = 8'haf;
memory[16'h0400] = 8'h2c;
memory[16'h0401] = 8'h03;
memory[16'h0402] = 8'h3c;
memory[16'h0403] = 8'h28;
memory[16'h0404] = 8'hd6;
memory[16'h0405] = 8'h04;
memory[16'h0406] = 8'h12;
memory[16'h0407] = 8'h7b;
memory[16'h0408] = 8'h15;
memory[16'h0409] = 8'hb0;
memory[16'h040a] = 8'he2;
memory[16'h040b] = 8'h44;
memory[16'h040c] = 8'h08;
memory[16'h040d] = 8'he2;
memory[16'h040e] = 8'h6b;
memory[16'h040f] = 8'h0d;
memory[16'h0410] = 8'h38;
memory[16'h0411] = 8'h09;
memory[16'h0412] = 8'h48;
memory[16'h0413] = 8'he0;
memory[16'h0414] = 8'h58;
memory[16'h0415] = 8'he1;
memory[16'h0416] = 8'hc2;
memory[16'h0417] = 8'h82;
memory[16'h0418] = 8'ha6;
memory[16'h0419] = 8'he8;
memory[16'h041a] = 8'hff;
memory[16'h041b] = 8'heb;
memory[16'h041c] = 8'h02;
memory[16'h041d] = 8'hcf;
memory[16'h041e] = 8'haf;
memory[16'h041f] = 8'ha0;
memory[16'h0420] = 8'he2;
memory[16'h0421] = 8'hc2;
memory[16'h0422] = 8'h72;
memory[16'h0423] = 8'hd6;
memory[16'h0424] = 8'h03;
memory[16'h0425] = 8'h91;
memory[16'h0426] = 8'heb;
memory[16'h0427] = 8'h14;
memory[16'h0428] = 8'h8a;
memory[16'h0429] = 8'hf5;
memory[16'h042a] = 8'hc2;
memory[16'h042b] = 8'h60;
memory[16'h042c] = 8'hd6;
memory[16'h042d] = 8'h03;
memory[16'h042e] = 8'he2;
memory[16'h042f] = 8'h7b;
memory[16'h0430] = 8'h0a;
memory[16'h0431] = 8'ha0;
memory[16'h0432] = 8'he2;
memory[16'h0433] = 8'hc2;
memory[16'h0434] = 8'h82;
memory[16'h0435] = 8'ha0;
memory[16'h0436] = 8'he2;
memory[16'h0437] = 8'hc2;
memory[16'h0438] = 8'h92;
memory[16'h0439] = 8'hdf;
memory[16'h043a] = 8'haf;
memory[16'h043b] = 8'h8e;
memory[16'h043c] = 8'h8e;
memory[16'h043d] = 8'h8e;
memory[16'h043e] = 8'h02;
memory[16'h043f] = 8'h38;
memory[16'h0440] = 8'h16;
memory[16'h0441] = 8'he2;
memory[16'h0442] = 8'h00;
memory[16'h0443] = 8'h08;
memory[16'h0444] = 8'he4;
memory[16'h0445] = 8'h18;
memory[16'h0446] = 8'he5;
memory[16'h0447] = 8'h8b;
memory[16'h0448] = 8'hcd;
memory[16'h0449] = 8'h80;
memory[16'h044a] = 8'he0;
memory[16'h044b] = 8'hd6;
memory[16'h044c] = 8'h04;
memory[16'h044d] = 8'h00;
memory[16'h044e] = 8'hc2;
memory[16'h044f] = 8'ha0;
memory[16'h0450] = 8'ha6;
memory[16'h0451] = 8'hea;
memory[16'h0452] = 8'h5b;
memory[16'h0453] = 8'heb;
memory[16'h0454] = 8'h1a;
memory[16'h0455] = 8'ha0;
memory[16'h0456] = 8'he0;
memory[16'h0457] = 8'h70;
memory[16'h0458] = 8'he8;
memory[16'h0459] = 8'h70;
memory[16'h045a] = 8'he9;
memory[16'h045b] = 8'hd6;
memory[16'h045c] = 8'h04;
memory[16'h045d] = 8'hc7;
memory[16'h045e] = 8'h50;
memory[16'h045f] = 8'he9;
memory[16'h0460] = 8'h50;
memory[16'h0461] = 8'he8;
memory[16'h0462] = 8'h7c;
memory[16'h0463] = 8'h5d;
memory[16'h0464] = 8'hd6;
memory[16'h0465] = 8'h03;
memory[16'h0466] = 8'h91;
memory[16'h0467] = 8'h6b;
memory[16'h0468] = 8'h06;
memory[16'h0469] = 8'h70;
memory[16'h046a] = 8'he3;
memory[16'h046b] = 8'h70;
memory[16'h046c] = 8'he2;
memory[16'h046d] = 8'h8b;
memory[16'h046e] = 8'he8;
memory[16'h046f] = 8'h48;
memory[16'h0470] = 8'he2;
memory[16'h0471] = 8'h58;
memory[16'h0472] = 8'he3;
memory[16'h0473] = 8'hd4;
memory[16'h0474] = 8'he8;
memory[16'h0475] = 8'h31;
memory[16'h0476] = 8'h10;
memory[16'h0477] = 8'hdf;
memory[16'h0478] = 8'haf;
memory[16'h0479] = 8'hd6;
memory[16'h047a] = 8'h03;
memory[16'h047b] = 8'hd9;
memory[16'h047c] = 8'hfb;
memory[16'h047d] = 8'h17;
memory[16'h047e] = 8'hc2;
memory[16'h047f] = 8'h70;
memory[16'h0480] = 8'hfe;
memory[16'h0481] = 8'hd6;
memory[16'h0482] = 8'h03;
memory[16'h0483] = 8'he2;
memory[16'h0484] = 8'h7b;
memory[16'h0485] = 8'hc3;
memory[16'h0486] = 8'h26;
memory[16'h0487] = 8'he6;
memory[16'h0488] = 8'h41;
memory[16'h0489] = 8'h90;
memory[16'h048a] = 8'he6;
memory[16'h048b] = 8'h06;
memory[16'h048c] = 8'he6;
memory[16'h048d] = 8'h20;
memory[16'h048e] = 8'he3;
memory[16'h048f] = 8'h26;
memory[16'h0490] = 8'h6e;
memory[16'h0491] = 8'he3;
memory[16'h0492] = 8'h36;
memory[16'h0493] = 8'hdf;
memory[16'h0494] = 8'haf;
memory[16'h0495] = 8'ha7;
memory[16'h0496] = 8'hef;
memory[16'h0497] = 8'h3b;
memory[16'h0498] = 8'h6b;
memory[16'h0499] = 8'h19;
memory[16'h049a] = 8'ha7;
memory[16'h049b] = 8'hef;
memory[16'h049c] = 8'h0d;
memory[16'h049d] = 8'h6b;
memory[16'h049e] = 8'h14;
memory[16'h049f] = 8'hfe;
memory[16'h04a0] = 8'hc3;
memory[16'h04a1] = 8'hf0;
memory[16'h04a2] = 8'h00;
memory[16'h04a3] = 8'hef;
memory[16'h04a4] = 8'hd6;
memory[16'h04a5] = 8'h03;
memory[16'h04a6] = 8'hf2;
memory[16'h04a7] = 8'hfe;
memory[16'h04a8] = 8'h7b;
memory[16'h04a9] = 8'hf6;
memory[16'h04aa] = 8'h80;
memory[16'h04ab] = 8'he0;
memory[16'h04ac] = 8'hd6;
memory[16'h04ad] = 8'h01;
memory[16'h04ae] = 8'hd9;
memory[16'h04af] = 8'h28;
memory[16'h04b0] = 8'he4;
memory[16'h04b1] = 8'h38;
memory[16'h04b2] = 8'he5;
memory[16'h04b3] = 8'haf;
memory[16'h04b4] = 8'h7c;
memory[16'h04b5] = 8'h28;
memory[16'h04b6] = 8'hd6;
memory[16'h04b7] = 8'h03;
memory[16'h04b8] = 8'h91;
memory[16'h04b9] = 8'heb;
memory[16'h04ba] = 8'hbe;
memory[16'h04bb] = 8'hd6;
memory[16'h04bc] = 8'h04;
memory[16'h04bd] = 8'hc7;
memory[16'h04be] = 8'hfb;
memory[16'h04bf] = 8'h06;
memory[16'h04c0] = 8'h7c;
memory[16'h04c1] = 8'h29;
memory[16'h04c2] = 8'hd6;
memory[16'h04c3] = 8'h03;
memory[16'h04c4] = 8'h91;
memory[16'h04c5] = 8'hef;
memory[16'h04c6] = 8'haf;
memory[16'h04c7] = 8'hd6;
memory[16'h04c8] = 8'h04;
memory[16'h04c9] = 8'hb4;
memory[16'h04ca] = 8'hfb;
memory[16'h04cb] = 8'h09;
memory[16'h04cc] = 8'hd6;
memory[16'h04cd] = 8'h03;
memory[16'h04ce] = 8'h91;
memory[16'h04cf] = 8'hd6;
memory[16'h04d0] = 8'h03;
memory[16'h04d1] = 8'h9a;
memory[16'h04d2] = 8'h6b;
memory[16'h04d3] = 8'h04;
memory[16'h04d4] = 8'hdf;
memory[16'h04d5] = 8'h80;
memory[16'h04d6] = 8'he0;
memory[16'h04d7] = 8'haf;
memory[16'h04d8] = 8'h70;
memory[16'h04d9] = 8'he8;
memory[16'h04da] = 8'h70;
memory[16'h04db] = 8'he9;
memory[16'h04dc] = 8'h70;
memory[16'h04dd] = 8'he2;
memory[16'h04de] = 8'h70;
memory[16'h04df] = 8'he3;
memory[16'h04e0] = 8'hd6;
memory[16'h04e1] = 8'h04;
memory[16'h04e2] = 8'hb4;
memory[16'h04e3] = 8'h48;
memory[16'h04e4] = 8'he2;
memory[16'h04e5] = 8'h58;
memory[16'h04e6] = 8'he3;
memory[16'h04e7] = 8'h50;
memory[16'h04e8] = 8'he3;
memory[16'h04e9] = 8'h50;
memory[16'h04ea] = 8'he2;
memory[16'h04eb] = 8'h50;
memory[16'h04ec] = 8'he9;
memory[16'h04ed] = 8'h50;
memory[16'h04ee] = 8'he8;
memory[16'h04ef] = 8'hd4;
memory[16'h04f0] = 8'he8;
memory[16'h04f1] = 8'h8b;
memory[16'h04f2] = 8'hd9;
memory[16'h04f3] = 8'hd6;
memory[16'h04f4] = 8'h03;
memory[16'h04f5] = 8'h91;
memory[16'h04f6] = 8'h26;
memory[16'h04f7] = 8'he6;
memory[16'h04f8] = 8'h41;
memory[16'h04f9] = 8'h02;
memory[16'h04fa] = 8'h66;
memory[16'h04fb] = 8'h8c;
memory[16'h04fc] = 8'h20;
memory[16'h04fd] = 8'h02;
memory[16'h04fe] = 8'h86;
memory[16'h04ff] = 8'haf;
memory[16'h0500] = 8'hc2;
memory[16'h0501] = 8'h40;
memory[16'h0502] = 8'h80;
memory[16'h0503] = 8'he0;
memory[16'h0504] = 8'h76;
memory[16'h0505] = 8'he4;
memory[16'h0506] = 8'h80;
memory[16'h0507] = 8'h6b;
memory[16'h0508] = 8'hf7;
memory[16'h0509] = 8'ha0;
memory[16'h050a] = 8'he0;
memory[16'h050b] = 8'h56;
memory[16'h050c] = 8'he4;
memory[16'h050d] = 8'h7f;
memory[16'h050e] = 8'ha4;
memory[16'h050f] = 8'h06;
memory[16'h0510] = 8'he0;
memory[16'h0511] = 8'heb;
memory[16'h0512] = 8'h06;
memory[16'h0513] = 8'ha4;
memory[16'h0514] = 8'h07;
memory[16'h0515] = 8'he1;
memory[16'h0516] = 8'hdf;
memory[16'h0517] = 8'h6b;
memory[16'h0518] = 8'h0f;
memory[16'h0519] = 8'h80;
memory[16'h051a] = 8'he0;
memory[16'h051b] = 8'hc2;
memory[16'h051c] = 8'h50;
memory[16'h051d] = 8'ha0;
memory[16'h051e] = 8'he0;
memory[16'h051f] = 8'ha6;
memory[16'h0520] = 8'he5;
memory[16'h0521] = 8'h0d;
memory[16'h0522] = 8'h6b;
memory[16'h0523] = 8'h04;
memory[16'h0524] = 8'h80;
memory[16'h0525] = 8'he0;
memory[16'h0526] = 8'h8b;
memory[16'h0527] = 8'hd8;
memory[16'h0528] = 8'ha0;
memory[16'h0529] = 8'he0;
memory[16'h052a] = 8'hc2;
memory[16'h052b] = 8'h50;
memory[16'h052c] = 8'h80;
memory[16'h052d] = 8'he0;
memory[16'h052e] = 8'haf;
memory[16'h052f] = 8'h7c;
memory[16'h0530] = 8'h22;
memory[16'h0531] = 8'hd6;
memory[16'h0532] = 8'h03;
memory[16'h0533] = 8'h91;
memory[16'h0534] = 8'heb;
memory[16'h0535] = 8'h0c;
memory[16'h0536] = 8'hd6;
memory[16'h0537] = 8'h03;
memory[16'h0538] = 8'h91;
memory[16'h0539] = 8'h6b;
memory[16'h053a] = 8'h09;
memory[16'h053b] = 8'h58;
memory[16'h053c] = 8'he6;
memory[16'h053d] = 8'hd6;
memory[16'h053e] = 8'h08;
memory[16'h053f] = 8'h18;
memory[16'h0540] = 8'h8b;
memory[16'h0541] = 8'hf4;
memory[16'h0542] = 8'h80;
memory[16'h0543] = 8'he0;
memory[16'h0544] = 8'haf;
memory[16'h0545] = 8'hd6;
memory[16'h0546] = 8'h04;
memory[16'h0547] = 8'hc7;
memory[16'h0548] = 8'hb0;
memory[16'h0549] = 8'hea;
memory[16'h054a] = 8'h9c;
memory[16'h054b] = 8'h02;
memory[16'h054c] = 8'h8c;
memory[16'h054d] = 8'h10;
memory[16'h054e] = 8'hc2;
memory[16'h054f] = 8'h60;
memory[16'h0550] = 8'ha6;
memory[16'h0551] = 8'he6;
memory[16'h0552] = 8'h3c;
memory[16'h0553] = 8'h6b;
memory[16'h0554] = 8'h0e;
memory[16'h0555] = 8'h90;
memory[16'h0556] = 8'he8;
memory[16'h0557] = 8'ha6;
memory[16'h0558] = 8'he6;
memory[16'h0559] = 8'h3e;
memory[16'h055a] = 8'h6b;
memory[16'h055b] = 8'h07;
memory[16'h055c] = 8'h90;
memory[16'h055d] = 8'he8;
memory[16'h055e] = 8'ha6;
memory[16'h055f] = 8'he6;
memory[16'h0560] = 8'h3d;
memory[16'h0561] = 8'heb;
memory[16'h0562] = 8'h06;
memory[16'h0563] = 8'h42;
memory[16'h0564] = 8'ha8;
memory[16'h0565] = 8'ha0;
memory[16'h0566] = 8'he0;
memory[16'h0567] = 8'h9a;
memory[16'h0568] = 8'he3;
memory[16'h0569] = 8'h70;
memory[16'h056a] = 8'hea;
memory[16'h056b] = 8'h70;
memory[16'h056c] = 8'he2;
memory[16'h056d] = 8'h70;
memory[16'h056e] = 8'he3;
memory[16'h056f] = 8'hd6;
memory[16'h0570] = 8'h04;
memory[16'h0571] = 8'hc7;
memory[16'h0572] = 8'h48;
memory[16'h0573] = 8'he2;
memory[16'h0574] = 8'h58;
memory[16'h0575] = 8'he3;
memory[16'h0576] = 8'h50;
memory[16'h0577] = 8'he3;
memory[16'h0578] = 8'h50;
memory[16'h0579] = 8'he2;
memory[16'h057a] = 8'hd6;
memory[16'h057b] = 8'h01;
memory[16'h057c] = 8'h41;
memory[16'h057d] = 8'h50;
memory[16'h057e] = 8'he8;
memory[16'h057f] = 8'h54;
memory[16'h0580] = 8'h0f;
memory[16'h0581] = 8'he8;
memory[16'h0582] = 8'haf;
memory[16'h0583] = 8'h7c;
memory[16'h0584] = 8'h3b;
memory[16'h0585] = 8'hd6;
memory[16'h0586] = 8'h03;
memory[16'h0587] = 8'h91;
memory[16'h0588] = 8'h6b;
memory[16'h0589] = 8'h06;
memory[16'h058a] = 8'ha6;
memory[16'h058b] = 8'he6;
memory[16'h058c] = 8'h0d;
memory[16'h058d] = 8'hdf;
memory[16'h058e] = 8'heb;
memory[16'h058f] = 8'hf5;
memory[16'h0590] = 8'h80;
memory[16'h0591] = 8'he0;
memory[16'h0592] = 8'haf;
memory[16'h0593] = 8'hd6;
memory[16'h0594] = 8'h05;
memory[16'h0595] = 8'h83;
memory[16'h0596] = 8'h7b;
memory[16'h0597] = 8'hfa;
memory[16'h0598] = 8'ha0;
memory[16'h0599] = 8'he0;
memory[16'h059a] = 8'h8b;
memory[16'h059b] = 8'hf7;
memory[16'h059c] = 8'hd6;
memory[16'h059d] = 8'h04;
memory[16'h059e] = 8'hf3;
memory[16'h059f] = 8'h70;
memory[16'h05a0] = 8'he8;
memory[16'h05a1] = 8'ha0;
memory[16'h05a2] = 8'he0;
memory[16'h05a3] = 8'hd6;
memory[16'h05a4] = 8'h04;
memory[16'h05a5] = 8'hc7;
memory[16'h05a6] = 8'h50;
memory[16'h05a7] = 8'he8;
memory[16'h05a8] = 8'hf3;
memory[16'h05a9] = 8'h82;
memory[16'h05aa] = 8'h8e;
memory[16'h05ab] = 8'hf3;
memory[16'h05ac] = 8'h83;
memory[16'h05ad] = 8'haf;
memory[16'h05ae] = 8'h09;
memory[16'h05af] = 8'h04;
memory[16'h05b0] = 8'h19;
memory[16'h05b1] = 8'h05;
memory[16'h05b2] = 8'h8b;
memory[16'h05b3] = 8'hcf;
memory[16'h05b4] = 8'h70;
memory[16'h05b5] = 8'h04;
memory[16'h05b6] = 8'h70;
memory[16'h05b7] = 8'h05;
memory[16'h05b8] = 8'h09;
memory[16'h05b9] = 8'h04;
memory[16'h05ba] = 8'h19;
memory[16'h05bb] = 8'h05;
memory[16'h05bc] = 8'hc2;
memory[16'h05bd] = 8'h60;
memory[16'h05be] = 8'ha6;
memory[16'h05bf] = 8'he6;
memory[16'h05c0] = 8'h5b;
memory[16'h05c1] = 8'heb;
memory[16'h05c2] = 8'h15;
memory[16'h05c3] = 8'ha0;
memory[16'h05c4] = 8'he0;
memory[16'h05c5] = 8'hb0;
memory[16'h05c6] = 8'he8;
memory[16'h05c7] = 8'h7c;
memory[16'h05c8] = 8'h5d;
memory[16'h05c9] = 8'ha0;
memory[16'h05ca] = 8'he0;
memory[16'h05cb] = 8'hd6;
memory[16'h05cc] = 8'h03;
memory[16'h05cd] = 8'h91;
memory[16'h05ce] = 8'h6b;
memory[16'h05cf] = 8'h06;
memory[16'h05d0] = 8'h70;
memory[16'h05d1] = 8'he8;
memory[16'h05d2] = 8'h70;
memory[16'h05d3] = 8'he8;
memory[16'h05d4] = 8'h8b;
memory[16'h05d5] = 8'hf3;
memory[16'h05d6] = 8'ha0;
memory[16'h05d7] = 8'he0;
memory[16'h05d8] = 8'hd6;
memory[16'h05d9] = 8'h04;
memory[16'h05da] = 8'h4b;
memory[16'h05db] = 8'h08;
memory[16'h05dc] = 8'h04;
memory[16'h05dd] = 8'h18;
memory[16'h05de] = 8'h05;
memory[16'h05df] = 8'h7c;
memory[16'h05e0] = 8'h5b;
memory[16'h05e1] = 8'hd6;
memory[16'h05e2] = 8'h03;
memory[16'h05e3] = 8'h91;
memory[16'h05e4] = 8'heb;
memory[16'h05e5] = 8'h18;
memory[16'h05e6] = 8'h7c;
memory[16'h05e7] = 8'h5d;
memory[16'h05e8] = 8'hd6;
memory[16'h05e9] = 8'h04;
memory[16'h05ea] = 8'hf3;
memory[16'h05eb] = 8'hd6;
memory[16'h05ec] = 8'h03;
memory[16'h05ed] = 8'h91;
memory[16'h05ee] = 8'h6b;
memory[16'h05ef] = 8'h0b;
memory[16'h05f0] = 8'h50;
memory[16'h05f1] = 8'hea;
memory[16'h05f2] = 8'hf3;
memory[16'h05f3] = 8'h8a;
memory[16'h05f4] = 8'h50;
memory[16'h05f5] = 8'hea;
memory[16'h05f6] = 8'h8e;
memory[16'h05f7] = 8'hf3;
memory[16'h05f8] = 8'h8a;
memory[16'h05f9] = 8'h8b;
memory[16'h05fa] = 8'hed;
memory[16'h05fb] = 8'hd6;
memory[16'h05fc] = 8'h05;
memory[16'h05fd] = 8'ha8;
memory[16'h05fe] = 8'h50;
memory[16'h05ff] = 8'h05;
memory[16'h0600] = 8'h50;
memory[16'h0601] = 8'h04;
memory[16'h0602] = 8'h8b;
memory[16'h0603] = 8'hae;
memory[16'h0604] = 8'hd6;
memory[16'h0605] = 8'h04;
memory[16'h0606] = 8'hc7;
memory[16'h0607] = 8'hd6;
memory[16'h0608] = 8'h05;
memory[16'h0609] = 8'h00;
memory[16'h060a] = 8'hd6;
memory[16'h060b] = 8'h01;
memory[16'h060c] = 8'h41;
memory[16'h060d] = 8'h76;
memory[16'h060e] = 8'h0f;
memory[16'h060f] = 8'h50;
memory[16'h0610] = 8'heb;
memory[16'h0611] = 8'h1f;
memory[16'h0612] = 8'hd6;
memory[16'h0613] = 8'h05;
memory[16'h0614] = 8'h93;
memory[16'h0615] = 8'ha0;
memory[16'h0616] = 8'he0;
memory[16'h0617] = 8'hc2;
memory[16'h0618] = 8'h40;
memory[16'h0619] = 8'ha0;
memory[16'h061a] = 8'he0;
memory[16'h061b] = 8'hc2;
memory[16'h061c] = 8'h50;
memory[16'h061d] = 8'h80;
memory[16'h061e] = 8'he0;
memory[16'h061f] = 8'h90;
memory[16'h0620] = 8'he4;
memory[16'h0621] = 8'hcf;
memory[16'h0622] = 8'hc0;
memory[16'h0623] = 8'he4;
memory[16'h0624] = 8'hfb;
memory[16'h0625] = 8'h08;
memory[16'h0626] = 8'hd6;
memory[16'h0627] = 8'h01;
memory[16'h0628] = 8'h41;
memory[16'h0629] = 8'h76;
memory[16'h062a] = 8'h0f;
memory[16'h062b] = 8'h50;
memory[16'h062c] = 8'h6b;
memory[16'h062d] = 8'he4;
memory[16'h062e] = 8'h80;
memory[16'h062f] = 8'he0;
memory[16'h0630] = 8'haf;
memory[16'h0631] = 8'hd6;
memory[16'h0632] = 8'h05;
memory[16'h0633] = 8'h00;
memory[16'h0634] = 8'hfb;
memory[16'h0635] = 8'h07;
memory[16'h0636] = 8'ha0;
memory[16'h0637] = 8'hfe;
memory[16'h0638] = 8'ha0;
memory[16'h0639] = 8'hfe;
memory[16'h063a] = 8'h8d;
memory[16'h063b] = 8'h07;
memory[16'h063c] = 8'h3e;
memory[16'h063d] = 8'hd6;
memory[16'h063e] = 8'h01;
memory[16'h063f] = 8'h41;
memory[16'h0640] = 8'h76;
memory[16'h0641] = 8'h0f;
memory[16'h0642] = 8'h60;
memory[16'h0643] = 8'heb;
memory[16'h0644] = 8'he9;
memory[16'h0645] = 8'h80;
memory[16'h0646] = 8'he0;
memory[16'h0647] = 8'h8b;
memory[16'h0648] = 8'he8;
memory[16'h0649] = 8'h56;
memory[16'h064a] = 8'h0f;
memory[16'h064b] = 8'hfe;
memory[16'h064c] = 8'hd6;
memory[16'h064d] = 8'h05;
memory[16'h064e] = 8'h45;
memory[16'h064f] = 8'heb;
memory[16'h0650] = 8'h05;
memory[16'h0651] = 8'h20;
memory[16'h0652] = 8'h0f;
memory[16'h0653] = 8'h8d;
memory[16'h0654] = 8'h05;
memory[16'h0655] = 8'h93;
memory[16'h0656] = 8'haf;
memory[16'h0657] = 8'h76;
memory[16'h0658] = 8'h0f;
memory[16'h0659] = 8'h01;
memory[16'h065a] = 8'h6d;
memory[16'h065b] = 8'h05;
memory[16'h065c] = 8'h93;
memory[16'h065d] = 8'h56;
memory[16'h065e] = 8'h0f;
memory[16'h065f] = 8'hfe;
memory[16'h0660] = 8'haf;
memory[16'h0661] = 8'ha6;
memory[16'h0662] = 8'h0e;
memory[16'h0663] = 8'h00;
memory[16'h0664] = 8'heb;
memory[16'h0665] = 8'h06;
memory[16'h0666] = 8'h46;
memory[16'h0667] = 8'h0e;
memory[16'h0668] = 8'h20;
memory[16'h0669] = 8'h8d;
memory[16'h066a] = 8'h01;
memory[16'h066b] = 8'h1b;
memory[16'h066c] = 8'h00;
memory[16'h066d] = 8'h0e;
memory[16'h066e] = 8'h50;
memory[16'h066f] = 8'he6;
memory[16'h0670] = 8'h50;
memory[16'h0671] = 8'he7;
memory[16'h0672] = 8'h50;
memory[16'h0673] = 8'he0;
memory[16'h0674] = 8'h50;
memory[16'h0675] = 8'he1;
memory[16'h0676] = 8'h56;
memory[16'h0677] = 8'h0f;
memory[16'h0678] = 8'hfe;
memory[16'h0679] = 8'h30;
memory[16'h067a] = 8'he6;
memory[16'h067b] = 8'h88;
memory[16'h067c] = 8'he0;
memory[16'h067d] = 8'h98;
memory[16'h067e] = 8'he1;
memory[16'h067f] = 8'hd6;
memory[16'h0680] = 8'h05;
memory[16'h0681] = 8'h83;
memory[16'h0682] = 8'h50;
memory[16'h0683] = 8'hea;
memory[16'h0684] = 8'h50;
memory[16'h0685] = 8'heb;
memory[16'h0686] = 8'h70;
memory[16'h0687] = 8'he1;
memory[16'h0688] = 8'h70;
memory[16'h0689] = 8'he0;
memory[16'h068a] = 8'h70;
memory[16'h068b] = 8'heb;
memory[16'h068c] = 8'h70;
memory[16'h068d] = 8'hea;
memory[16'h068e] = 8'h08;
memory[16'h068f] = 8'he8;
memory[16'h0690] = 8'h18;
memory[16'h0691] = 8'he9;
memory[16'h0692] = 8'h20;
memory[16'h0693] = 8'h0e;
memory[16'h0694] = 8'h76;
memory[16'h0695] = 8'h0e;
memory[16'h0696] = 8'h10;
memory[16'h0697] = 8'h6d;
memory[16'h0698] = 8'h06;
memory[16'h0699] = 8'h04;
memory[16'h069a] = 8'hd6;
memory[16'h069b] = 8'h05;
memory[16'h069c] = 8'h83;
memory[16'h069d] = 8'h8b;
memory[16'h069e] = 8'hca;
memory[16'h069f] = 8'hd6;
memory[16'h06a0] = 8'h04;
memory[16'h06a1] = 8'hc7;
memory[16'h06a2] = 8'h68;
memory[16'h06a3] = 8'he2;
memory[16'h06a4] = 8'h42;
memory[16'h06a5] = 8'h63;
memory[16'h06a6] = 8'h6b;
memory[16'h06a7] = 8'h10;
memory[16'h06a8] = 8'h40;
memory[16'h06a9] = 8'he6;
memory[16'h06aa] = 8'h6c;
memory[16'h06ab] = 8'h00;
memory[16'h06ac] = 8'h7c;
memory[16'h06ad] = 8'hb4;
memory[16'h06ae] = 8'h80;
memory[16'h06af] = 8'he6;
memory[16'h06b0] = 8'hed;
memory[16'h06b1] = 8'h06;
memory[16'h06b2] = 8'hae;
memory[16'h06b3] = 8'h80;
memory[16'h06b4] = 8'he2;
memory[16'h06b5] = 8'hed;
memory[16'h06b6] = 8'h06;
memory[16'h06b7] = 8'ha8;
memory[16'h06b8] = 8'haf;
memory[16'h06b9] = 8'hd6;
memory[16'h06ba] = 8'h04;
memory[16'h06bb] = 8'hc7;
memory[16'h06bc] = 8'hd4;
memory[16'h06bd] = 8'he2;
memory[16'h06be] = 8'h31;
memory[16'h06bf] = 8'h10;
memory[16'h06c0] = 8'haf;
memory[16'h06c1] = 8'h46;
memory[16'h06c2] = 8'h0f;
memory[16'h06c3] = 8'h08;
memory[16'h06c4] = 8'haf;
memory[16'h06c5] = 8'h46;
memory[16'h06c6] = 8'h0f;
memory[16'h06c7] = 8'h02;
memory[16'h06c8] = 8'haf;
memory[16'h06c9] = 8'hb0;
memory[16'h06ca] = 8'h04;
memory[16'h06cb] = 8'hb0;
memory[16'h06cc] = 8'h05;
memory[16'h06cd] = 8'haf;
memory[16'h06ce] = 8'hd6;
memory[16'h06cf] = 8'h05;
memory[16'h06d0] = 8'h2f;
memory[16'h06d1] = 8'hd6;
memory[16'h06d2] = 8'h04;
memory[16'h06d3] = 8'hc7;
memory[16'h06d4] = 8'hfb;
memory[16'h06d5] = 8'h22;
memory[16'h06d6] = 8'hd6;
memory[16'h06d7] = 8'h01;
memory[16'h06d8] = 8'h5e;
memory[16'h06d9] = 8'hac;
memory[16'h06da] = 8'h05;
memory[16'h06db] = 8'h8b;
memory[16'h06dc] = 8'h0d;
memory[16'h06dd] = 8'hd6;
memory[16'h06de] = 8'h05;
memory[16'h06df] = 8'h2f;
memory[16'h06e0] = 8'hd6;
memory[16'h06e1] = 8'h04;
memory[16'h06e2] = 8'hc7;
memory[16'h06e3] = 8'hfb;
memory[16'h06e4] = 8'h13;
memory[16'h06e5] = 8'hd6;
memory[16'h06e6] = 8'h01;
memory[16'h06e7] = 8'h82;
memory[16'h06e8] = 8'hac;
memory[16'h06e9] = 8'h06;
memory[16'h06ea] = 8'hbc;
memory[16'h06eb] = 8'h14;
memory[16'h06ec] = 8'h70;
memory[16'h06ed] = 8'he5;
memory[16'h06ee] = 8'he3;
memory[16'h06ef] = 8'h5b;
memory[16'h06f0] = 8'hbe;
memory[16'h06f1] = 8'hd6;
memory[16'h06f2] = 8'h08;
memory[16'h06f3] = 8'h18;
memory[16'h06f4] = 8'h50;
memory[16'h06f5] = 8'he5;
memory[16'h06f6] = 8'haa;
memory[16'h06f7] = 8'hf4;
memory[16'h06f8] = 8'hc2;
memory[16'h06f9] = 8'h60;
memory[16'h06fa] = 8'ha6;
memory[16'h06fb] = 8'he6;
memory[16'h06fc] = 8'h2c;
memory[16'h06fd] = 8'heb;
memory[16'h06fe] = 8'h11;
memory[16'h06ff] = 8'ha0;
memory[16'h0700] = 8'he0;
memory[16'h0701] = 8'hc2;
memory[16'h0702] = 8'h60;
memory[16'h0703] = 8'ha6;
memory[16'h0704] = 8'he6;
memory[16'h0705] = 8'h3b;
memory[16'h0706] = 8'h6b;
memory[16'h0707] = 8'h07;
memory[16'h0708] = 8'ha6;
memory[16'h0709] = 8'he6;
memory[16'h070a] = 8'h0d;
memory[16'h070b] = 8'h6b;
memory[16'h070c] = 8'h02;
memory[16'h070d] = 8'h80;
memory[16'h070e] = 8'he0;
memory[16'h070f] = 8'haf;
memory[16'h0710] = 8'h5c;
memory[16'h0711] = 8'h0d;
memory[16'h0712] = 8'h8d;
memory[16'h0713] = 8'h08;
memory[16'h0714] = 8'h18;
memory[16'h0715] = 8'hd6;
memory[16'h0716] = 8'h05;
memory[16'h0717] = 8'h2f;
memory[16'h0718] = 8'hd6;
memory[16'h0719] = 8'h02;
memory[16'h071a] = 8'he9;
memory[16'h071b] = 8'hd6;
memory[16'h071c] = 8'h04;
memory[16'h071d] = 8'hf3;
memory[16'h071e] = 8'h8d;
memory[16'h071f] = 8'h05;
memory[16'h0720] = 8'ha8;
memory[16'h0721] = 8'he6;
memory[16'h0722] = 8'h0f;
memory[16'h0723] = 8'h04;
memory[16'h0724] = 8'h8b;
memory[16'h0725] = 8'h10;
memory[16'h0726] = 8'he6;
memory[16'h0727] = 8'h0f;
memory[16'h0728] = 8'h08;
memory[16'h0729] = 8'h8b;
memory[16'h072a] = 8'h0b;
memory[16'h072b] = 8'hb0;
memory[16'h072c] = 8'h0f;
memory[16'h072d] = 8'hb0;
memory[16'h072e] = 8'h0e;
memory[16'h072f] = 8'h08;
memory[16'h0730] = 8'h06;
memory[16'h0731] = 8'h18;
memory[16'h0732] = 8'h07;
memory[16'h0733] = 8'hd6;
memory[16'h0734] = 8'h06;
memory[16'h0735] = 8'hc9;
memory[16'h0736] = 8'h31;
memory[16'h0737] = 8'h10;
memory[16'h0738] = 8'h50;
memory[16'h0739] = 8'h0a;
memory[16'h073a] = 8'h50;
memory[16'h073b] = 8'h0b;
memory[16'h073c] = 8'h8b;
memory[16'h073d] = 8'h0a;
memory[16'h073e] = 8'h76;
memory[16'h073f] = 8'h0f;
memory[16'h0740] = 8'h0a;
memory[16'h0741] = 8'heb;
memory[16'h0742] = 8'h0a;
memory[16'h0743] = 8'h66;
memory[16'h0744] = 8'h0f;
memory[16'h0745] = 8'h84;
memory[16'h0746] = 8'h6b;
memory[16'h0747] = 8'h05;
memory[16'h0748] = 8'hc2;
memory[16'h0749] = 8'h60;
memory[16'h074a] = 8'h6e;
memory[16'h074b] = 8'h6a;
memory[16'h074c] = 8'h02;
memory[16'h074d] = 8'h30;
memory[16'h074e] = 8'h0a;
memory[16'h074f] = 8'ha4;
memory[16'h0750] = 8'he0;
memory[16'h0751] = 8'h06;
memory[16'h0752] = 8'heb;
memory[16'h0753] = 8'h05;
memory[16'h0754] = 8'ha4;
memory[16'h0755] = 8'he1;
memory[16'h0756] = 8'h07;
memory[16'h0757] = 8'h6b;
memory[16'h0758] = 8'h2c;
memory[16'h0759] = 8'h68;
memory[16'h075a] = 8'h04;
memory[16'h075b] = 8'h44;
memory[16'h075c] = 8'h05;
memory[16'h075d] = 8'he6;
memory[16'h075e] = 8'h6b;
memory[16'h075f] = 8'h25;
memory[16'h0760] = 8'h70;
memory[16'h0761] = 8'he1;
memory[16'h0762] = 8'h70;
memory[16'h0763] = 8'he0;
memory[16'h0764] = 8'h08;
memory[16'h0765] = 8'h04;
memory[16'h0766] = 8'h18;
memory[16'h0767] = 8'h05;
memory[16'h0768] = 8'hd6;
memory[16'h0769] = 8'h05;
memory[16'h076a] = 8'h45;
memory[16'h076b] = 8'h6b;
memory[16'h076c] = 8'h14;
memory[16'h076d] = 8'hd6;
memory[16'h076e] = 8'h06;
memory[16'h076f] = 8'hc9;
memory[16'h0770] = 8'h50;
memory[16'h0771] = 8'he6;
memory[16'h0772] = 8'h50;
memory[16'h0773] = 8'he7;
memory[16'h0774] = 8'h80;
memory[16'h0775] = 8'he6;
memory[16'h0776] = 8'h70;
memory[16'h0777] = 8'he7;
memory[16'h0778] = 8'h70;
memory[16'h0779] = 8'he6;
memory[16'h077a] = 8'ha0;
memory[16'h077b] = 8'he0;
memory[16'h077c] = 8'hd6;
memory[16'h077d] = 8'h06;
memory[16'h077e] = 8'h92;
memory[16'h077f] = 8'h8b;
memory[16'h0780] = 8'h38;
memory[16'h0781] = 8'h50;
memory[16'h0782] = 8'he0;
memory[16'h0783] = 8'h50;
memory[16'h0784] = 8'he1;
memory[16'h0785] = 8'ha0;
memory[16'h0786] = 8'he0;
memory[16'h0787] = 8'ha0;
memory[16'h0788] = 8'he0;
memory[16'h0789] = 8'hc2;
memory[16'h078a] = 8'h30;
memory[16'h078b] = 8'ha0;
memory[16'h078c] = 8'he0;
memory[16'h078d] = 8'ha6;
memory[16'h078e] = 8'he3;
memory[16'h078f] = 8'h3e;
memory[16'h0790] = 8'h6b;
memory[16'h0791] = 8'h03;
memory[16'h0792] = 8'h56;
memory[16'h0793] = 8'h0f;
memory[16'h0794] = 8'hfe;
memory[16'h0795] = 8'h6c;
memory[16'h0796] = 8'h07;
memory[16'h0797] = 8'h7c;
memory[16'h0798] = 8'hc8;
memory[16'h0799] = 8'hb0;
memory[16'h079a] = 8'he2;
memory[16'h079b] = 8'hc2;
memory[16'h079c] = 8'h86;
memory[16'h079d] = 8'ha2;
memory[16'h079e] = 8'h83;
memory[16'h079f] = 8'h6b;
memory[16'h07a0] = 8'h05;
memory[16'h07a1] = 8'ha0;
memory[16'h07a2] = 8'he6;
memory[16'h07a3] = 8'h2e;
memory[16'h07a4] = 8'h8b;
memory[16'h07a5] = 8'hf5;
memory[16'h07a6] = 8'h02;
memory[16'h07a7] = 8'h22;
memory[16'h07a8] = 8'h6c;
memory[16'h07a9] = 8'h07;
memory[16'h07aa] = 8'h7c;
memory[16'h07ab] = 8'hd9;
memory[16'h07ac] = 8'h02;
memory[16'h07ad] = 8'h72;
memory[16'h07ae] = 8'h16;
memory[16'h07af] = 8'he6;
memory[16'h07b0] = 8'h00;
memory[16'h07b1] = 8'h2c;
memory[16'h07b2] = 8'h0c;
memory[16'h07b3] = 8'hc3;
memory[16'h07b4] = 8'h26;
memory[16'h07b5] = 8'hc3;
memory[16'h07b6] = 8'h26;
memory[16'h07b7] = 8'hd4;
memory[16'h07b8] = 8'h0c;
memory[16'h07b9] = 8'h7c;
memory[16'h07ba] = 8'h0d;
memory[16'h07bb] = 8'hd6;
memory[16'h07bc] = 8'h03;
memory[16'h07bd] = 8'h91;
memory[16'h07be] = 8'h6d;
memory[16'h07bf] = 8'h07;
memory[16'h07c0] = 8'h3e;
memory[16'h07c1] = 8'ha6;
memory[16'h07c2] = 8'he6;
memory[16'h07c3] = 8'h3b;
memory[16'h07c4] = 8'h6b;
memory[16'h07c5] = 8'hc3;
memory[16'h07c6] = 8'h8b;
memory[16'h07c7] = 8'hef;
memory[16'h07c8] = 8'h4c;
memory[16'h07c9] = 8'h4f;
memory[16'h07ca] = 8'h47;
memory[16'h07cb] = 8'h46;
memory[16'h07cc] = 8'h3e;
memory[16'h07cd] = 8'h52;
memory[16'h07ce] = 8'h53;
memory[16'h07cf] = 8'h57;
memory[16'h07d0] = 8'h4d;
memory[16'h07d1] = 8'h43;
memory[16'h07d2] = 8'h54;
memory[16'h07d3] = 8'h45;
memory[16'h07d4] = 8'h21;
memory[16'h07d5] = 8'h2f;
memory[16'h07d6] = 8'h50;
memory[16'h07d7] = 8'h48;
memory[16'h07d8] = 8'h49;
memory[16'h07d9] = 8'h05;
memory[16'h07da] = 8'h9c;
memory[16'h07db] = 8'h05;
memory[16'h07dc] = 8'hb4;
memory[16'h07dd] = 8'h06;
memory[16'h07de] = 8'h04;
memory[16'h07df] = 8'h06;
memory[16'h07e0] = 8'h49;
memory[16'h07e1] = 8'h06;
memory[16'h07e2] = 8'h57;
memory[16'h07e3] = 8'h06;
memory[16'h07e4] = 8'h61;
memory[16'h07e5] = 8'h06;
memory[16'h07e6] = 8'h7b;
memory[16'h07e7] = 8'h06;
memory[16'h07e8] = 8'h9f;
memory[16'h07e9] = 8'h05;
memory[16'h07ea] = 8'h83;
memory[16'h07eb] = 8'h06;
memory[16'h07ec] = 8'hb9;
memory[16'h07ed] = 8'h06;
memory[16'h07ee] = 8'hc1;
memory[16'h07ef] = 8'h06;
memory[16'h07f0] = 8'hc5;
memory[16'h07f1] = 8'h05;
memory[16'h07f2] = 8'hae;
memory[16'h07f3] = 8'h06;
memory[16'h07f4] = 8'hc9;
memory[16'h07f5] = 8'h06;
memory[16'h07f6] = 8'hdd;
memory[16'h07f7] = 8'h06;
memory[16'h07f8] = 8'hce;
memory[16'h07f9] = 8'h07;
memory[16'h07fa] = 8'h15;
memory[16'h07fb] = 8'hff;
memory[16'h07fc] = 8'hff;
memory[16'h07fd] = 8'h8d;
memory[16'h07fe] = 8'h07;
memory[16'h07ff] = 8'h2b;
memory[16'h0800] = 8'h8d;
memory[16'h0801] = 8'he0;
memory[16'h0802] = 8'h00;
memory[16'h0803] = 8'h8d;
memory[16'h0804] = 8'he0;
memory[16'h0805] = 8'h03;
memory[16'h0806] = 8'h8d;
memory[16'h0807] = 8'he0;
memory[16'h0808] = 8'h06;
memory[16'h0809] = 8'h8d;
memory[16'h080a] = 8'he0;
memory[16'h080b] = 8'h09;
memory[16'h080c] = 8'h8d;
memory[16'h080d] = 8'h0a;
memory[16'h080e] = 8'hda;
memory[16'h080f] = 8'h8d;
memory[16'h0810] = 8'he0;
memory[16'h0811] = 8'h0f;
memory[16'h0812] = 8'h8d;
memory[16'h0813] = 8'h08;
memory[16'h0814] = 8'hff;
memory[16'h0815] = 8'h8d;
memory[16'h0816] = 8'h08;
memory[16'h0817] = 8'h1d;
memory[16'h0818] = 8'he4;
memory[16'h0819] = 8'h15;
memory[16'h081a] = 8'h5a;
memory[16'h081b] = 8'h8b;
memory[16'h081c] = 8'h0a;
memory[16'h081d] = 8'hd6;
memory[16'h081e] = 8'h08;
memory[16'h081f] = 8'h24;
memory[16'h0820] = 8'he4;
memory[16'h0821] = 8'h5a;
memory[16'h0822] = 8'h13;
memory[16'h0823] = 8'haf;
memory[16'h0824] = 8'hd6;
memory[16'h0825] = 8'h0c;
memory[16'h0826] = 8'h1d;
memory[16'h0827] = 8'ha6;
memory[16'h0828] = 8'h5a;
memory[16'h0829] = 8'h7f;
memory[16'h082a] = 8'h6b;
memory[16'h082b] = 8'h3f;
memory[16'h082c] = 8'ha6;
memory[16'h082d] = 8'h5a;
memory[16'h082e] = 8'h20;
memory[16'h082f] = 8'hfb;
memory[16'h0830] = 8'h41;
memory[16'h0831] = 8'ha6;
memory[16'h0832] = 8'h5a;
memory[16'h0833] = 8'h1b;
memory[16'h0834] = 8'h6b;
memory[16'h0835] = 8'h3f;
memory[16'h0836] = 8'he6;
memory[16'h0837] = 8'h5c;
memory[16'h0838] = 8'hf0;
memory[16'h0839] = 8'ha6;
memory[16'h083a] = 8'h5a;
memory[16'h083b] = 8'h1a;
memory[16'h083c] = 8'h6b;
memory[16'h083d] = 8'h3a;
memory[16'h083e] = 8'he6;
memory[16'h083f] = 8'h5c;
memory[16'h0840] = 8'h10;
memory[16'h0841] = 8'ha6;
memory[16'h0842] = 8'h5a;
memory[16'h0843] = 8'h0a;
memory[16'h0844] = 8'h6b;
memory[16'h0845] = 8'h32;
memory[16'h0846] = 8'he6;
memory[16'h0847] = 8'h5c;
memory[16'h0848] = 8'hff;
memory[16'h0849] = 8'ha6;
memory[16'h084a] = 8'h5a;
memory[16'h084b] = 8'h0b;
memory[16'h084c] = 8'h6b;
memory[16'h084d] = 8'h2a;
memory[16'h084e] = 8'ha6;
memory[16'h084f] = 8'h5a;
memory[16'h0850] = 8'h08;
memory[16'h0851] = 8'heb;
memory[16'h0852] = 8'h0d;
memory[16'h0853] = 8'hd6;
memory[16'h0854] = 8'h08;
memory[16'h0855] = 8'h78;
memory[16'h0856] = 8'he6;
memory[16'h0857] = 8'h5a;
memory[16'h0858] = 8'h20;
memory[16'h0859] = 8'hd6;
memory[16'h085a] = 8'h0b;
memory[16'h085b] = 8'h95;
memory[16'h085c] = 8'he6;
memory[16'h085d] = 8'h5a;
memory[16'h085e] = 8'h08;
memory[16'h085f] = 8'haf;
memory[16'h0860] = 8'ha6;
memory[16'h0861] = 8'h5a;
memory[16'h0862] = 8'h0d;
memory[16'h0863] = 8'heb;
memory[16'h0864] = 8'h07;
memory[16'h0865] = 8'hd6;
memory[16'h0866] = 8'h0a;
memory[16'h0867] = 8'hd4;
memory[16'h0868] = 8'he6;
memory[16'h0869] = 8'h5a;
memory[16'h086a] = 8'h0d;
memory[16'h086b] = 8'haf;
memory[16'h086c] = 8'ha6;
memory[16'h086d] = 8'h5a;
memory[16'h086e] = 8'h0c;
memory[16'h086f] = 8'h6b;
memory[16'h0870] = 8'h6c;
memory[16'h0871] = 8'haf;
memory[16'h0872] = 8'hd6;
memory[16'h0873] = 8'h0b;
memory[16'h0874] = 8'h95;
memory[16'h0875] = 8'he6;
memory[16'h0876] = 8'h5c;
memory[16'h0877] = 8'h01;
memory[16'h0878] = 8'h04;
memory[16'h0879] = 8'h5c;
memory[16'h087a] = 8'h5b;
memory[16'h087b] = 8'h4b;
memory[16'h087c] = 8'h1c;
memory[16'h087d] = 8'h5b;
memory[16'h087e] = 8'h7d;
memory[16'h087f] = 8'he4;
memory[16'h0880] = 8'h5c;
memory[16'h0881] = 8'h60;
memory[16'h0882] = 8'he4;
memory[16'h0883] = 8'h5b;
memory[16'h0884] = 8'h5c;
memory[16'h0885] = 8'h56;
memory[16'h0886] = 8'h5c;
memory[16'h0887] = 8'h0f;
memory[16'h0888] = 8'ha6;
memory[16'h0889] = 8'h5c;
memory[16'h088a] = 8'h0d;
memory[16'h088b] = 8'h7b;
memory[16'h088c] = 8'h4f;
memory[16'h088d] = 8'h90;
memory[16'h088e] = 8'h60;
memory[16'h088f] = 8'hfb;
memory[16'h0890] = 8'h03;
memory[16'h0891] = 8'h26;
memory[16'h0892] = 8'h5b;
memory[16'h0893] = 8'h06;
memory[16'h0894] = 8'h06;
memory[16'h0895] = 8'h5b;
memory[16'h0896] = 8'h03;
memory[16'h0897] = 8'hcb;
memory[16'h0898] = 8'h43;
memory[16'h0899] = 8'h70;
memory[16'h089a] = 8'hfd;
memory[16'h089b] = 8'h31;
memory[16'h089c] = 8'h60;
memory[16'h089d] = 8'h0c;
memory[16'h089e] = 8'hfd;
memory[16'h089f] = 8'h1c;
memory[16'h08a0] = 8'h00;
memory[16'h08a1] = 8'h2c;
memory[16'h08a2] = 8'hfd;
memory[16'h08a3] = 8'h3c;
memory[16'h08a4] = 8'h10;
memory[16'h08a5] = 8'h4c;
memory[16'h08a6] = 8'h70;
memory[16'h08a7] = 8'h82;
memory[16'h08a8] = 8'h52;
memory[16'h08a9] = 8'h92;
memory[16'h08aa] = 8'h50;
memory[16'h08ab] = 8'h1e;
memory[16'h08ac] = 8'h3e;
memory[16'h08ad] = 8'h4a;
memory[16'h08ae] = 8'hf8;
memory[16'h08af] = 8'h4c;
memory[16'h08b0] = 8'h10;
memory[16'h08b1] = 8'h5c;
memory[16'h08b2] = 8'h20;
memory[16'h08b3] = 8'h92;
memory[16'h08b4] = 8'h50;
memory[16'h08b5] = 8'h1e;
memory[16'h08b6] = 8'h4a;
memory[16'h08b7] = 8'hfb;
memory[16'h08b8] = 8'h1c;
memory[16'h08b9] = 8'h38;
memory[16'h08ba] = 8'h2e;
memory[16'h08bb] = 8'h0e;
memory[16'h08bc] = 8'h3c;
memory[16'h08bd] = 8'h70;
memory[16'h08be] = 8'h39;
memory[16'h08bf] = 8'h5b;
memory[16'h08c0] = 8'h82;
memory[16'h08c1] = 8'h52;
memory[16'h08c2] = 8'h92;
memory[16'h08c3] = 8'h50;
memory[16'h08c4] = 8'ha0;
memory[16'h08c5] = 8'he0;
memory[16'h08c6] = 8'ha0;
memory[16'h08c7] = 8'he2;
memory[16'h08c8] = 8'ha6;
memory[16'h08c9] = 8'he3;
memory[16'h08ca] = 8'hf0;
memory[16'h08cb] = 8'h7b;
memory[16'h08cc] = 8'hf3;
memory[16'h08cd] = 8'h5c;
memory[16'h08ce] = 8'hff;
memory[16'h08cf] = 8'ha2;
memory[16'h08d0] = 8'h25;
memory[16'h08d1] = 8'h7b;
memory[16'h08d2] = 8'hed;
memory[16'h08d3] = 8'h4c;
memory[16'h08d4] = 8'h38;
memory[16'h08d5] = 8'h92;
memory[16'h08d6] = 8'h50;
memory[16'h08d7] = 8'h1e;
memory[16'h08d8] = 8'h4a;
memory[16'h08d9] = 8'hfb;
memory[16'h08da] = 8'h50;
memory[16'h08db] = 8'hfd;
memory[16'h08dc] = 8'haf;
memory[16'h08dd] = 8'h70;
memory[16'h08de] = 8'hfd;
memory[16'h08df] = 8'h31;
memory[16'h08e0] = 8'h60;
memory[16'h08e1] = 8'h4c;
memory[16'h08e2] = 8'hfd;
memory[16'h08e3] = 8'h5c;
memory[16'h08e4] = 8'h80;
memory[16'h08e5] = 8'h3c;
memory[16'h08e6] = 8'h20;
memory[16'h08e7] = 8'h2c;
memory[16'h08e8] = 8'h80;
memory[16'h08e9] = 8'h00;
memory[16'h08ea] = 8'he5;
memory[16'h08eb] = 8'h92;
memory[16'h08ec] = 8'h34;
memory[16'h08ed] = 8'h2a;
memory[16'h08ee] = 8'hfa;
memory[16'h08ef] = 8'h2c;
memory[16'h08f0] = 8'h02;
memory[16'h08f1] = 8'h3c;
memory[16'h08f2] = 8'hff;
memory[16'h08f3] = 8'h4e;
memory[16'h08f4] = 8'h92;
memory[16'h08f5] = 8'h34;
memory[16'h08f6] = 8'h5a;
memory[16'h08f7] = 8'hfc;
memory[16'h08f8] = 8'h2a;
memory[16'h08f9] = 8'hf9;
memory[16'h08fa] = 8'h50;
memory[16'h08fb] = 8'hfd;
memory[16'h08fc] = 8'hb0;
memory[16'h08fd] = 8'h5b;
memory[16'h08fe] = 8'haf;
memory[16'h08ff] = 8'h31;
memory[16'h0900] = 8'hf0;
memory[16'h0901] = 8'hfc;
memory[16'h0902] = 8'h00;
memory[16'h0903] = 8'hec;
memory[16'h0904] = 8'hfe;
memory[16'h0905] = 8'hbc;
memory[16'h0906] = 8'h10;
memory[16'h0907] = 8'h9c;
memory[16'h0908] = 8'h08;
memory[16'h0909] = 8'h8c;
memory[16'h090a] = 8'h92;
memory[16'h090b] = 8'h5c;
memory[16'h090c] = 8'h05;
memory[16'h090d] = 8'h4c;
memory[16'h090e] = 8'h40;
memory[16'h090f] = 8'h1c;
memory[16'h0910] = 8'h03;
memory[16'h0911] = 8'he6;
memory[16'h0912] = 8'h06;
memory[16'h0913] = 8'he0;
memory[16'h0914] = 8'hb0;
memory[16'h0915] = 8'h07;
memory[16'h0916] = 8'hb0;
memory[16'h0917] = 8'h08;
memory[16'h0918] = 8'hb0;
memory[16'h0919] = 8'h6d;
memory[16'h091a] = 8'hd6;
memory[16'h091b] = 8'h08;
memory[16'h091c] = 8'hdd;
memory[16'h091d] = 8'h9f;
memory[16'h091e] = 8'he6;
memory[16'h091f] = 8'h58;
memory[16'h0920] = 8'h14;
memory[16'h0921] = 8'hd6;
memory[16'h0922] = 8'h0b;
memory[16'h0923] = 8'hf2;
memory[16'h0924] = 8'h31;
memory[16'h0925] = 8'h10;
memory[16'h0926] = 8'he6;
memory[16'h0927] = 8'h5a;
memory[16'h0928] = 8'h4b;
memory[16'h0929] = 8'hd6;
memory[16'h092a] = 8'h0b;
memory[16'h092b] = 8'h95;
memory[16'h092c] = 8'hd6;
memory[16'h092d] = 8'h08;
memory[16'h092e] = 8'h24;
memory[16'h092f] = 8'h68;
memory[16'h0930] = 8'h5a;
memory[16'h0931] = 8'hfc;
memory[16'h0932] = 8'h16;
memory[16'h0933] = 8'hd6;
memory[16'h0934] = 8'h03;
memory[16'h0935] = 8'hd9;
memory[16'h0936] = 8'hfb;
memory[16'h0937] = 8'h15;
memory[16'h0938] = 8'h26;
memory[16'h0939] = 8'he6;
memory[16'h093a] = 8'h31;
memory[16'h093b] = 8'h02;
memory[16'h093c] = 8'h66;
memory[16'h093d] = 8'he3;
memory[16'h093e] = 8'h26;
memory[16'h093f] = 8'h6e;
memory[16'h0940] = 8'he3;
memory[16'h0941] = 8'h36;
memory[16'h0942] = 8'he6;
memory[16'h0943] = 8'h5a;
memory[16'h0944] = 8'h3d;
memory[16'h0945] = 8'hd6;
memory[16'h0946] = 8'h08;
memory[16'h0947] = 8'h72;
memory[16'h0948] = 8'hd6;
memory[16'h0949] = 8'h0e;
memory[16'h094a] = 8'h92;
memory[16'h094b] = 8'h8b;
memory[16'h094c] = 8'hd7;
memory[16'h094d] = 8'ha6;
memory[16'h094e] = 8'he6;
memory[16'h094f] = 8'h2a;
memory[16'h0950] = 8'heb;
memory[16'h0951] = 8'h0a;
memory[16'h0952] = 8'h76;
memory[16'h0953] = 8'h0f;
memory[16'h0954] = 8'h08;
memory[16'h0955] = 8'h6b;
memory[16'h0956] = 8'h36;
memory[16'h0957] = 8'h56;
memory[16'h0958] = 8'h0f;
memory[16'h0959] = 8'hf7;
memory[16'h095a] = 8'h8b;
memory[16'h095b] = 8'h1c;
memory[16'h095c] = 8'he6;
memory[16'h095d] = 8'h0f;
memory[16'h095e] = 8'h04;
memory[16'h095f] = 8'hb0;
memory[16'h0960] = 8'h0e;
memory[16'h0961] = 8'h08;
memory[16'h0962] = 8'h06;
memory[16'h0963] = 8'h18;
memory[16'h0964] = 8'h07;
memory[16'h0965] = 8'ha6;
memory[16'h0966] = 8'he6;
memory[16'h0967] = 8'h08;
memory[16'h0968] = 8'heb;
memory[16'h0969] = 8'h06;
memory[16'h096a] = 8'h4c;
memory[16'h096b] = 8'h00;
memory[16'h096c] = 8'h92;
memory[16'h096d] = 8'h40;
memory[16'h096e] = 8'h8b;
memory[16'h096f] = 8'hb4;
memory[16'h0970] = 8'ha6;
memory[16'h0971] = 8'he6;
memory[16'h0972] = 8'h2b;
memory[16'h0973] = 8'heb;
memory[16'h0974] = 8'h36;
memory[16'h0975] = 8'hd6;
memory[16'h0976] = 8'h06;
memory[16'h0977] = 8'hc9;
memory[16'h0978] = 8'hd6;
memory[16'h0979] = 8'h07;
memory[16'h097a] = 8'h38;
memory[16'h097b] = 8'hd6;
memory[16'h097c] = 8'h0a;
memory[16'h097d] = 8'hd4;
memory[16'h097e] = 8'he6;
memory[16'h097f] = 8'h58;
memory[16'h0980] = 8'h0c;
memory[16'h0981] = 8'h76;
memory[16'h0982] = 8'h0f;
memory[16'h0983] = 8'h02;
memory[16'h0984] = 8'heb;
memory[16'h0985] = 8'h0c;
memory[16'h0986] = 8'h00;
memory[16'h0987] = 8'h58;
memory[16'h0988] = 8'h76;
memory[16'h0989] = 8'h0f;
memory[16'h098a] = 8'h08;
memory[16'h098b] = 8'heb;
memory[16'h098c] = 8'h05;
memory[16'h098d] = 8'hd6;
memory[16'h098e] = 8'h0e;
memory[16'h098f] = 8'h80;
memory[16'h0990] = 8'h8b;
memory[16'h0991] = 8'h92;
memory[16'h0992] = 8'hd6;
memory[16'h0993] = 8'h0b;
memory[16'h0994] = 8'hf2;
memory[16'h0995] = 8'h70;
memory[16'h0996] = 8'he0;
memory[16'h0997] = 8'h70;
memory[16'h0998] = 8'he1;
memory[16'h0999] = 8'h80;
memory[16'h099a] = 8'he0;
memory[16'h099b] = 8'hd6;
memory[16'h099c] = 8'h05;
memory[16'h099d] = 8'h00;
memory[16'h099e] = 8'h28;
memory[16'h099f] = 8'he4;
memory[16'h09a0] = 8'h38;
memory[16'h09a1] = 8'he5;
memory[16'h09a2] = 8'hd6;
memory[16'h09a3] = 8'h0e;
memory[16'h09a4] = 8'h92;
memory[16'h09a5] = 8'h50;
memory[16'h09a6] = 8'he1;
memory[16'h09a7] = 8'h50;
memory[16'h09a8] = 8'he0;
memory[16'h09a9] = 8'h8b;
memory[16'h09aa] = 8'he5;
memory[16'h09ab] = 8'ha6;
memory[16'h09ac] = 8'he6;
memory[16'h09ad] = 8'h2d;
memory[16'h09ae] = 8'he6;
memory[16'h09af] = 8'h6e;
memory[16'h09b0] = 8'h0c;
memory[16'h09b1] = 8'heb;
memory[16'h09b2] = 8'h26;
memory[16'h09b3] = 8'he6;
memory[16'h09b4] = 8'h6f;
memory[16'h09b5] = 8'he6;
memory[16'h09b6] = 8'h82;
memory[16'h09b7] = 8'h20;
memory[16'h09b8] = 8'h42;
memory[16'h09b9] = 8'h22;
memory[16'h09ba] = 8'h6b;
memory[16'h09bb] = 8'hd4;
memory[16'h09bc] = 8'ha0;
memory[16'h09bd] = 8'he0;
memory[16'h09be] = 8'h82;
memory[16'h09bf] = 8'h30;
memory[16'h09c0] = 8'h56;
memory[16'h09c1] = 8'he2;
memory[16'h09c2] = 8'h7f;
memory[16'h09c3] = 8'hd6;
memory[16'h09c4] = 8'h0a;
memory[16'h09c5] = 8'ha3;
memory[16'h09c6] = 8'hd6;
memory[16'h09c7] = 8'h0d;
memory[16'h09c8] = 8'hcc;
memory[16'h09c9] = 8'hfb;
memory[16'h09ca] = 8'hc2;
memory[16'h09cb] = 8'hb0;
memory[16'h09cc] = 8'h6d;
memory[16'h09cd] = 8'hd6;
memory[16'h09ce] = 8'h0c;
memory[16'h09cf] = 8'h1d;
memory[16'h09d0] = 8'ha6;
memory[16'h09d1] = 8'h5a;
memory[16'h09d2] = 8'h2d;
memory[16'h09d3] = 8'heb;
memory[16'h09d4] = 8'hbb;
memory[16'h09d5] = 8'ha0;
memory[16'h09d6] = 8'he0;
memory[16'h09d7] = 8'h8b;
memory[16'h09d8] = 8'hdd;
memory[16'h09d9] = 8'hd6;
memory[16'h09da] = 8'h03;
memory[16'h09db] = 8'he7;
memory[16'h09dc] = 8'hfb;
memory[16'h09dd] = 8'h5a;
memory[16'h09de] = 8'h38;
memory[16'h09df] = 8'he6;
memory[16'h09e0] = 8'hd6;
memory[16'h09e1] = 8'h02;
memory[16'h09e2] = 8'hf4;
memory[16'h09e3] = 8'hfc;
memory[16'h09e4] = 8'h16;
memory[16'h09e5] = 8'h8c;
memory[16'h09e6] = 8'h80;
memory[16'h09e7] = 8'h42;
memory[16'h09e8] = 8'h84;
memory[16'h09e9] = 8'h98;
memory[16'h09ea] = 8'he5;
memory[16'h09eb] = 8'h42;
memory[16'h09ec] = 8'h95;
memory[16'h09ed] = 8'heb;
memory[16'h09ee] = 8'h01;
memory[16'h09ef] = 8'h9e;
memory[16'h09f0] = 8'h82;
memory[16'h09f1] = 8'h20;
memory[16'h09f2] = 8'h42;
memory[16'h09f3] = 8'h22;
memory[16'h09f4] = 8'h6b;
memory[16'h09f5] = 8'h1d;
memory[16'h09f6] = 8'h56;
memory[16'h09f7] = 8'he2;
memory[16'h09f8] = 8'h7f;
memory[16'h09f9] = 8'ha0;
memory[16'h09fa] = 8'he0;
memory[16'h09fb] = 8'h82;
memory[16'h09fc] = 8'h30;
memory[16'h09fd] = 8'hd6;
memory[16'h09fe] = 8'h01;
memory[16'h09ff] = 8'h41;
memory[16'h0a00] = 8'h76;
memory[16'h0a01] = 8'h0f;
memory[16'h0a02] = 8'h40;
memory[16'h0a03] = 8'heb;
memory[16'h0a04] = 8'h2e;
memory[16'h0a05] = 8'h76;
memory[16'h0a06] = 8'h0f;
memory[16'h0a07] = 8'h20;
memory[16'h0a08] = 8'heb;
memory[16'h0a09] = 8'h07;
memory[16'h0a0a] = 8'hd6;
memory[16'h0a0b] = 8'h05;
memory[16'h0a0c] = 8'h93;
memory[16'h0a0d] = 8'ha0;
memory[16'h0a0e] = 8'he0;
memory[16'h0a0f] = 8'h8b;
memory[16'h0a10] = 8'hdf;
memory[16'h0a11] = 8'h80;
memory[16'h0a12] = 8'he0;
memory[16'h0a13] = 8'he6;
memory[16'h0a14] = 8'h6f;
memory[16'h0a15] = 8'hd7;
memory[16'h0a16] = 8'h68;
memory[16'h0a17] = 8'he8;
memory[16'h0a18] = 8'hd6;
memory[16'h0a19] = 8'h0c;
memory[16'h0a1a] = 8'ha4;
memory[16'h0a1b] = 8'h68;
memory[16'h0a1c] = 8'he9;
memory[16'h0a1d] = 8'hd6;
memory[16'h0a1e] = 8'h0d;
memory[16'h0a1f] = 8'hcc;
memory[16'h0a20] = 8'h7b;
memory[16'h0a21] = 8'h0b;
memory[16'h0a22] = 8'hd6;
memory[16'h0a23] = 8'h0a;
memory[16'h0a24] = 8'h81;
memory[16'h0a25] = 8'h6e;
memory[16'h0a26] = 8'h5b;
memory[16'h0a27] = 8'h08;
memory[16'h0a28] = 8'hd6;
memory[16'h0a29] = 8'h0e;
memory[16'h0a2a] = 8'h80;
memory[16'h0a2b] = 8'h8b;
memory[16'h0a2c] = 8'h03;
memory[16'h0a2d] = 8'hd6;
memory[16'h0a2e] = 8'h0c;
memory[16'h0a2f] = 8'ha4;
memory[16'h0a30] = 8'h8d;
memory[16'h0a31] = 8'h09;
memory[16'h0a32] = 8'h24;
memory[16'h0a33] = 8'hd6;
memory[16'h0a34] = 8'h0a;
memory[16'h0a35] = 8'h81;
memory[16'h0a36] = 8'h8b;
memory[16'h0a37] = 8'hdb;
memory[16'h0a38] = 8'h8f;
memory[16'h0a39] = 8'he6;
memory[16'h0a3a] = 8'hf5;
memory[16'h0a3b] = 8'h21;
memory[16'h0a3c] = 8'he6;
memory[16'h0a3d] = 8'hf4;
memory[16'h0a3e] = 8'h0d;
memory[16'h0a3f] = 8'he6;
memory[16'h0a40] = 8'hf1;
memory[16'h0a41] = 8'h43;
memory[16'h0a42] = 8'he6;
memory[16'h0a43] = 8'hf7;
memory[16'h0a44] = 8'h48;
memory[16'h0a45] = 8'he6;
memory[16'h0a46] = 8'hf0;
memory[16'h0a47] = 8'hff;
memory[16'h0a48] = 8'hb0;
memory[16'h0a49] = 8'hfa;
memory[16'h0a4a] = 8'ha6;
memory[16'h0a4b] = 8'he6;
memory[16'h0a4c] = 8'h5f;
memory[16'h0a4d] = 8'heb;
memory[16'h0a4e] = 8'h14;
memory[16'h0a4f] = 8'h76;
memory[16'h0a50] = 8'hfa;
memory[16'h0a51] = 8'h08;
memory[16'h0a52] = 8'h6b;
memory[16'h0a53] = 8'hfb;
memory[16'h0a54] = 8'hb0;
memory[16'h0a55] = 8'hfa;
memory[16'h0a56] = 8'h68;
memory[16'h0a57] = 8'hf0;
memory[16'h0a58] = 8'h92;
memory[16'h0a59] = 8'h60;
memory[16'h0a5a] = 8'ha0;
memory[16'h0a5b] = 8'he0;
memory[16'h0a5c] = 8'h42;
memory[16'h0a5d] = 8'h66;
memory[16'h0a5e] = 8'heb;
memory[16'h0a5f] = 8'hef;
memory[16'h0a60] = 8'h8d;
memory[16'h0a61] = 8'h00;
memory[16'h0a62] = 8'h20;
memory[16'h0a63] = 8'ha6;
memory[16'h0a64] = 8'he6;
memory[16'h0a65] = 8'h40;
memory[16'h0a66] = 8'heb;
memory[16'h0a67] = 8'hf8;
memory[16'h0a68] = 8'h2c;
memory[16'h0a69] = 8'h14;
memory[16'h0a6a] = 8'hd6;
memory[16'h0a6b] = 8'h06;
memory[16'h0a6c] = 8'haa;
memory[16'h0a6d] = 8'h6e;
memory[16'h0a6e] = 8'h76;
memory[16'h0a6f] = 8'hfa;
memory[16'h0a70] = 8'h10;
memory[16'h0a71] = 8'h6b;
memory[16'h0a72] = 8'hfb;
memory[16'h0a73] = 8'hb0;
memory[16'h0a74] = 8'hfa;
memory[16'h0a75] = 8'h42;
memory[16'h0a76] = 8'h66;
memory[16'h0a77] = 8'h6b;
memory[16'h0a78] = 8'he7;
memory[16'h0a79] = 8'h82;
memory[16'h0a7a] = 8'h60;
memory[16'h0a7b] = 8'h69;
memory[16'h0a7c] = 8'hf0;
memory[16'h0a7d] = 8'ha0;
memory[16'h0a7e] = 8'he0;
memory[16'h0a7f] = 8'h8b;
memory[16'h0a80] = 8'hed;
memory[16'h0a81] = 8'hd6;
memory[16'h0a82] = 8'h05;
memory[16'h0a83] = 8'h00;
memory[16'h0a84] = 8'h28;
memory[16'h0a85] = 8'he0;
memory[16'h0a86] = 8'h38;
memory[16'h0a87] = 8'he1;
memory[16'h0a88] = 8'h48;
memory[16'h0a89] = 8'he0;
memory[16'h0a8a] = 8'h58;
memory[16'h0a8b] = 8'he1;
memory[16'h0a8c] = 8'ha0;
memory[16'h0a8d] = 8'he4;
memory[16'h0a8e] = 8'ha0;
memory[16'h0a8f] = 8'he4;
memory[16'h0a90] = 8'h82;
memory[16'h0a91] = 8'h74;
memory[16'h0a92] = 8'h90;
memory[16'h0a93] = 8'he7;
memory[16'h0a94] = 8'hbb;
memory[16'h0a95] = 8'hf8;
memory[16'h0a96] = 8'h82;
memory[16'h0a97] = 8'h74;
memory[16'h0a98] = 8'h92;
memory[16'h0a99] = 8'h72;
memory[16'h0a9a] = 8'ha0;
memory[16'h0a9b] = 8'he2;
memory[16'h0a9c] = 8'ha0;
memory[16'h0a9d] = 8'he4;
memory[16'h0a9e] = 8'h42;
memory[16'h0a9f] = 8'h77;
memory[16'h0aa0] = 8'heb;
memory[16'h0aa1] = 8'hf4;
memory[16'h0aa2] = 8'haf;
memory[16'h0aa3] = 8'hd6;
memory[16'h0aa4] = 8'h01;
memory[16'h0aa5] = 8'h82;
memory[16'h0aa6] = 8'ha6;
memory[16'h0aa7] = 8'he4;
memory[16'h0aa8] = 8'h20;
memory[16'h0aa9] = 8'h6b;
memory[16'h0aaa] = 8'h03;
memory[16'h0aab] = 8'hd6;
memory[16'h0aac] = 8'h0a;
memory[16'h0aad] = 8'hbd;
memory[16'h0aae] = 8'hbc;
memory[16'h0aaf] = 8'h15;
memory[16'h0ab0] = 8'he3;
memory[16'h0ab1] = 8'h4b;
memory[16'h0ab2] = 8'ha6;
memory[16'h0ab3] = 8'he4;
memory[16'h0ab4] = 8'h30;
memory[16'h0ab5] = 8'heb;
memory[16'h0ab6] = 8'h0b;
memory[16'h0ab7] = 8'hbe;
memory[16'h0ab8] = 8'ha6;
memory[16'h0ab9] = 8'heb;
memory[16'h0aba] = 8'h1a;
memory[16'h0abb] = 8'h7b;
memory[16'h0abc] = 8'hf3;
memory[16'h0abd] = 8'h49;
memory[16'h0abe] = 8'h5a;
memory[16'h0abf] = 8'h8d;
memory[16'h0ac0] = 8'h08;
memory[16'h0ac1] = 8'h72;
memory[16'h0ac2] = 8'hd6;
memory[16'h0ac3] = 8'h0a;
memory[16'h0ac4] = 8'hbd;
memory[16'h0ac5] = 8'hbe;
memory[16'h0ac6] = 8'he3;
memory[16'h0ac7] = 8'h4b;
memory[16'h0ac8] = 8'ha6;
memory[16'h0ac9] = 8'heb;
memory[16'h0aca] = 8'h1a;
memory[16'h0acb] = 8'h7b;
memory[16'h0acc] = 8'hf5;
memory[16'h0acd] = 8'haf;
memory[16'h0ace] = 8'he6;
memory[16'h0acf] = 8'h5a;
memory[16'h0ad0] = 8'h20;
memory[16'h0ad1] = 8'hd6;
memory[16'h0ad2] = 8'h08;
memory[16'h0ad3] = 8'h72;
memory[16'h0ad4] = 8'h76;
memory[16'h0ad5] = 8'h5b;
memory[16'h0ad6] = 8'h0f;
memory[16'h0ad7] = 8'heb;
memory[16'h0ad8] = 8'hf5;
memory[16'h0ad9] = 8'haf;
memory[16'h0ada] = 8'h70;
memory[16'h0adb] = 8'hfd;
memory[16'h0adc] = 8'h31;
memory[16'h0add] = 8'h50;
memory[16'h0ade] = 8'h4a;
memory[16'h0adf] = 8'h5e;
memory[16'h0ae0] = 8'h68;
memory[16'h0ae1] = 8'hfe;
memory[16'h0ae2] = 8'h78;
memory[16'h0ae3] = 8'hff;
memory[16'h0ae4] = 8'he6;
memory[16'h0ae5] = 8'hfe;
memory[16'h0ae6] = 8'hfe;
memory[16'h0ae7] = 8'hb0;
memory[16'h0ae8] = 8'hff;
memory[16'h0ae9] = 8'h4c;
memory[16'h0aea] = 8'h40;
memory[16'h0aeb] = 8'hf0;
memory[16'h0aec] = 8'h80;
memory[16'h0aed] = 8'h46;
memory[16'h0aee] = 8'h03;
memory[16'h0aef] = 8'h80;
memory[16'h0af0] = 8'h56;
memory[16'h0af1] = 8'h03;
memory[16'h0af2] = 8'h7f;
memory[16'h0af3] = 8'h76;
memory[16'h0af4] = 8'h6d;
memory[16'h0af5] = 8'h80;
memory[16'h0af6] = 8'h6b;
memory[16'h0af7] = 8'h05;
memory[16'h0af8] = 8'hb6;
memory[16'h0af9] = 8'h03;
memory[16'h0afa] = 8'h40;
memory[16'h0afb] = 8'h8b;
memory[16'h0afc] = 8'h05;
memory[16'h0afd] = 8'h56;
memory[16'h0afe] = 8'h03;
memory[16'h0aff] = 8'h3f;
memory[16'h0b00] = 8'h0b;
memory[16'h0b01] = 8'hfe;
memory[16'h0b02] = 8'h0b;
memory[16'h0b03] = 8'hfe;
memory[16'h0b04] = 8'hff;
memory[16'h0b05] = 8'h50;
memory[16'h0b06] = 8'h80;
memory[16'h0b07] = 8'hff;
memory[16'h0b08] = 8'h50;
memory[16'h0b09] = 8'h80;
memory[16'h0b0a] = 8'hff;
memory[16'h0b0b] = 8'h50;
memory[16'h0b0c] = 8'h80;
memory[16'h0b0d] = 8'hff;
memory[16'h0b0e] = 8'h50;
memory[16'h0b0f] = 8'h80;
memory[16'h0b10] = 8'hff;
memory[16'h0b11] = 8'h50;
memory[16'h0b12] = 8'h80;
memory[16'h0b13] = 8'hff;
memory[16'h0b14] = 8'h50;
memory[16'h0b15] = 8'h80;
memory[16'h0b16] = 8'hff;
memory[16'h0b17] = 8'h50;
memory[16'h0b18] = 8'h80;
memory[16'h0b19] = 8'hff;
memory[16'h0b1a] = 8'h50;
memory[16'h0b1b] = 8'h80;
memory[16'h0b1c] = 8'h5e;
memory[16'h0b1d] = 8'h6b;
memory[16'h0b1e] = 8'h08;
memory[16'h0b1f] = 8'h26;
memory[16'h0b20] = 8'hff;
memory[16'h0b21] = 8'h08;
memory[16'h0b22] = 8'h36;
memory[16'h0b23] = 8'hfe;
memory[16'h0b24] = 8'h00;
memory[16'h0b25] = 8'h8b;
memory[16'h0b26] = 8'hc4;
memory[16'h0b27] = 8'h5c;
memory[16'h0b28] = 8'hfd;
memory[16'h0b29] = 8'hff;
memory[16'h0b2a] = 8'hff;
memory[16'h0b2b] = 8'h4a;
memory[16'h0b2c] = 8'hbe;
memory[16'h0b2d] = 8'h56;
memory[16'h0b2e] = 8'hfa;
memory[16'h0b2f] = 8'hef;
memory[16'h0b30] = 8'h46;
memory[16'h0b31] = 8'h03;
memory[16'h0b32] = 8'h80;
memory[16'h0b33] = 8'h56;
memory[16'h0b34] = 8'h03;
memory[16'h0b35] = 8'h7f;
memory[16'h0b36] = 8'h69;
memory[16'h0b37] = 8'hfe;
memory[16'h0b38] = 8'h79;
memory[16'h0b39] = 8'hff;
memory[16'h0b3a] = 8'h4c;
memory[16'h0b3b] = 8'h78;
memory[16'h0b3c] = 8'h8b;
memory[16'h0b3d] = 8'h1c;
memory[16'h0b3e] = 8'ha6;
memory[16'h0b3f] = 8'he4;
memory[16'h0b40] = 8'h20;
memory[16'h0b41] = 8'h7b;
memory[16'h0b42] = 8'h0d;
memory[16'h0b43] = 8'ha6;
memory[16'h0b44] = 8'he4;
memory[16'h0b45] = 8'h25;
memory[16'h0b46] = 8'hfb;
memory[16'h0b47] = 8'h0c;
memory[16'h0b48] = 8'h56;
memory[16'h0b49] = 8'h03;
memory[16'h0b4a] = 8'h7f;
memory[16'h0b4b] = 8'h46;
memory[16'h0b4c] = 8'h03;
memory[16'h0b4d] = 8'h80;
memory[16'h0b4e] = 8'h8b;
memory[16'h0b4f] = 8'h0a;
memory[16'h0b50] = 8'ha0;
memory[16'h0b51] = 8'h56;
memory[16'h0b52] = 8'h80;
memory[16'h0b53] = 8'h56;
memory[16'h0b54] = 8'h46;
memory[16'h0b55] = 8'h03;
memory[16'h0b56] = 8'h80;
memory[16'h0b57] = 8'h56;
memory[16'h0b58] = 8'h03;
memory[16'h0b59] = 8'h7f;
memory[16'h0b5a] = 8'h50;
memory[16'h0b5b] = 8'hfd;
memory[16'h0b5c] = 8'hbf;
memory[16'h0b5d] = 8'h18;
memory[16'h0b5e] = 8'he2;
memory[16'h0b5f] = 8'h02;
memory[16'h0b60] = 8'h12;
memory[16'h0b61] = 8'h02;
memory[16'h0b62] = 8'h12;
memory[16'h0b63] = 8'h06;
memory[16'h0b64] = 8'he1;
memory[16'h0b65] = 8'he0;
memory[16'h0b66] = 8'h0c;
memory[16'h0b67] = 8'h0f;
memory[16'h0b68] = 8'haf;
memory[16'h0b69] = 8'h58;
memory[16'h0b6a] = 8'h5b;
memory[16'h0b6b] = 8'h56;
memory[16'h0b6c] = 8'he5;
memory[16'h0b6d] = 8'h0f;
memory[16'h0b6e] = 8'h38;
memory[16'h0b6f] = 8'he5;
memory[16'h0b70] = 8'h90;
memory[16'h0b71] = 8'he5;
memory[16'h0b72] = 8'h90;
memory[16'h0b73] = 8'he5;
memory[16'h0b74] = 8'h02;
memory[16'h0b75] = 8'h35;
memory[16'h0b76] = 8'h58;
memory[16'h0b77] = 8'he3;
memory[16'h0b78] = 8'h56;
memory[16'h0b79] = 8'he3;
memory[16'h0b7a] = 8'h07;
memory[16'h0b7b] = 8'h56;
memory[16'h0b7c] = 8'he5;
memory[16'h0b7d] = 8'h38;
memory[16'h0b7e] = 8'h90;
memory[16'h0b7f] = 8'he5;
memory[16'h0b80] = 8'hf0;
memory[16'h0b81] = 8'he5;
memory[16'h0b82] = 8'h68;
memory[16'h0b83] = 8'h5b;
memory[16'h0b84] = 8'hf0;
memory[16'h0b85] = 8'he6;
memory[16'h0b86] = 8'h4c;
memory[16'h0b87] = 8'hfe;
memory[16'h0b88] = 8'h56;
memory[16'h0b89] = 8'he6;
memory[16'h0b8a] = 8'h07;
memory[16'h0b8b] = 8'h6e;
memory[16'h0b8c] = 8'h06;
memory[16'h0b8d] = 8'he5;
memory[16'h0b8e] = 8'h38;
memory[16'h0b8f] = 8'h16;
memory[16'h0b90] = 8'he4;
memory[16'h0b91] = 8'h00;
memory[16'h0b92] = 8'h6a;
memory[16'h0b93] = 8'hf8;
memory[16'h0b94] = 8'haf;
memory[16'h0b95] = 8'h70;
memory[16'h0b96] = 8'hfd;
memory[16'h0b97] = 8'h31;
memory[16'h0b98] = 8'h60;
memory[16'h0b99] = 8'h0c;
memory[16'h0b9a] = 8'hfd;
memory[16'h0b9b] = 8'h18;
memory[16'h0b9c] = 8'h5b;
memory[16'h0b9d] = 8'h28;
memory[16'h0b9e] = 8'h5a;
memory[16'h0b9f] = 8'h92;
memory[16'h0ba0] = 8'h20;
memory[16'h0ba1] = 8'hd6;
memory[16'h0ba2] = 8'h0b;
memory[16'h0ba3] = 8'h5d;
memory[16'h0ba4] = 8'h2c;
memory[16'h0ba5] = 8'h03;
memory[16'h0ba6] = 8'hd6;
memory[16'h0ba7] = 8'h0b;
memory[16'h0ba8] = 8'h69;
memory[16'h0ba9] = 8'hc2;
memory[16'h0baa] = 8'h60;
memory[16'h0bab] = 8'hd6;
memory[16'h0bac] = 8'h0b;
memory[16'h0bad] = 8'hbb;
memory[16'h0bae] = 8'hc2;
memory[16'h0baf] = 8'h60;
memory[16'h0bb0] = 8'hf0;
memory[16'h0bb1] = 8'he6;
memory[16'h0bb2] = 8'hd6;
memory[16'h0bb3] = 8'h0b;
memory[16'h0bb4] = 8'hbb;
memory[16'h0bb5] = 8'h1e;
memory[16'h0bb6] = 8'h2a;
memory[16'h0bb7] = 8'hf1;
memory[16'h0bb8] = 8'h50;
memory[16'h0bb9] = 8'hfd;
memory[16'h0bba] = 8'haf;
memory[16'h0bbb] = 8'h82;
memory[16'h0bbc] = 8'h74;
memory[16'h0bbd] = 8'ha0;
memory[16'h0bbe] = 8'he4;
memory[16'h0bbf] = 8'h82;
memory[16'h0bc0] = 8'h84;
memory[16'h0bc1] = 8'h42;
memory[16'h0bc2] = 8'h33;
memory[16'h0bc3] = 8'h6b;
memory[16'h0bc4] = 8'h0a;
memory[16'h0bc5] = 8'ha8;
memory[16'h0bc6] = 8'he3;
memory[16'h0bc7] = 8'h90;
memory[16'h0bc8] = 8'he8;
memory[16'h0bc9] = 8'h10;
memory[16'h0bca] = 8'he7;
memory[16'h0bcb] = 8'h10;
memory[16'h0bcc] = 8'he9;
memory[16'h0bcd] = 8'haa;
memory[16'h0bce] = 8'hf8;
memory[16'h0bcf] = 8'h56;
memory[16'h0bd0] = 8'he7;
memory[16'h0bd1] = 8'h0f;
memory[16'h0bd2] = 8'h56;
memory[16'h0bd3] = 8'he6;
memory[16'h0bd4] = 8'hf0;
memory[16'h0bd5] = 8'h42;
memory[16'h0bd6] = 8'h76;
memory[16'h0bd7] = 8'h42;
memory[16'h0bd8] = 8'h33;
memory[16'h0bd9] = 8'h6b;
memory[16'h0bda] = 8'h0a;
memory[16'h0bdb] = 8'ha8;
memory[16'h0bdc] = 8'he3;
memory[16'h0bdd] = 8'he0;
memory[16'h0bde] = 8'he9;
memory[16'h0bdf] = 8'hc0;
memory[16'h0be0] = 8'he7;
memory[16'h0be1] = 8'hc0;
memory[16'h0be2] = 8'he8;
memory[16'h0be3] = 8'haa;
memory[16'h0be4] = 8'hf8;
memory[16'h0be5] = 8'h92;
memory[16'h0be6] = 8'h84;
memory[16'h0be7] = 8'h80;
memory[16'h0be8] = 8'he4;
memory[16'h0be9] = 8'h92;
memory[16'h0bea] = 8'h74;
memory[16'h0beb] = 8'h06;
memory[16'h0bec] = 8'he5;
memory[16'h0bed] = 8'h08;
memory[16'h0bee] = 8'h16;
memory[16'h0bef] = 8'he4;
memory[16'h0bf0] = 8'h00;
memory[16'h0bf1] = 8'haf;
memory[16'h0bf2] = 8'h70;
memory[16'h0bf3] = 8'hfd;
memory[16'h0bf4] = 8'h31;
memory[16'h0bf5] = 8'h50;
memory[16'h0bf6] = 8'hec;
memory[16'h0bf7] = 8'h0e;
memory[16'h0bf8] = 8'hfc;
memory[16'h0bf9] = 8'h98;
memory[16'h0bfa] = 8'h9c;
memory[16'h0bfb] = 8'h5a;
memory[16'h0bfc] = 8'hc3;
memory[16'h0bfd] = 8'h9e;
memory[16'h0bfe] = 8'h76;
memory[16'h0bff] = 8'hea;
memory[16'h0c00] = 8'h80;
memory[16'h0c01] = 8'h6b;
memory[16'h0c02] = 8'hf7;
memory[16'h0c03] = 8'h00;
memory[16'h0c04] = 8'he8;
memory[16'h0c05] = 8'heb;
memory[16'h0c06] = 8'hf3;
memory[16'h0c07] = 8'h56;
memory[16'h0c08] = 8'hea;
memory[16'h0c09] = 8'h7f;
memory[16'h0c0a] = 8'hd6;
memory[16'h0c0b] = 8'h08;
memory[16'h0c0c] = 8'h27;
memory[16'h0c0d] = 8'h9c;
memory[16'h0c0e] = 8'h5a;
memory[16'h0c0f] = 8'hc3;
memory[16'h0c10] = 8'h9e;
memory[16'h0c11] = 8'h76;
memory[16'h0c12] = 8'hea;
memory[16'h0c13] = 8'h80;
memory[16'h0c14] = 8'h6b;
memory[16'h0c15] = 8'hf4;
memory[16'h0c16] = 8'hac;
memory[16'h0c17] = 8'h20;
memory[16'h0c18] = 8'h50;
memory[16'h0c19] = 8'hfd;
memory[16'h0c1a] = 8'h8d;
memory[16'h0c1b] = 8'h08;
memory[16'h0c1c] = 8'h72;
memory[16'h0c1d] = 8'ha6;
memory[16'h0c1e] = 8'h54;
memory[16'h0c1f] = 8'h77;
memory[16'h0c20] = 8'heb;
memory[16'h0c21] = 8'hfb;
memory[16'h0c22] = 8'h70;
memory[16'h0c23] = 8'hfd;
memory[16'h0c24] = 8'h31;
memory[16'h0c25] = 8'h60;
memory[16'h0c26] = 8'h2c;
memory[16'h0c27] = 8'h05;
memory[16'h0c28] = 8'hd6;
memory[16'h0c29] = 8'h0b;
memory[16'h0c2a] = 8'h69;
memory[16'h0c2b] = 8'h6c;
memory[16'h0c2c] = 8'h00;
memory[16'h0c2d] = 8'hd6;
memory[16'h0c2e] = 8'h0b;
memory[16'h0c2f] = 8'hbb;
memory[16'h0c30] = 8'h2a;
memory[16'h0c31] = 8'hf9;
memory[16'h0c32] = 8'h0c;
memory[16'h0c33] = 8'hfd;
memory[16'h0c34] = 8'h18;
memory[16'h0c35] = 8'h5b;
memory[16'h0c36] = 8'h82;
memory[16'h0c37] = 8'h20;
memory[16'h0c38] = 8'h29;
memory[16'h0c39] = 8'h5a;
memory[16'h0c3a] = 8'h50;
memory[16'h0c3b] = 8'hfd;
memory[16'h0c3c] = 8'ha6;
memory[16'h0c3d] = 8'h54;
memory[16'h0c3e] = 8'h77;
memory[16'h0c3f] = 8'heb;
memory[16'h0c40] = 8'hfb;
memory[16'h0c41] = 8'hd6;
memory[16'h0c42] = 8'h0b;
memory[16'h0c43] = 8'h95;
memory[16'h0c44] = 8'hd6;
memory[16'h0c45] = 8'h0c;
memory[16'h0c46] = 8'h56;
memory[16'h0c47] = 8'h76;
memory[16'h0c48] = 8'h6d;
memory[16'h0c49] = 8'h7f;
memory[16'h0c4a] = 8'h6b;
memory[16'h0c4b] = 8'hd1;
memory[16'h0c4c] = 8'he4;
memory[16'h0c4d] = 8'h6d;
memory[16'h0c4e] = 8'h5a;
memory[16'h0c4f] = 8'h56;
memory[16'h0c50] = 8'h6d;
memory[16'h0c51] = 8'h80;
memory[16'h0c52] = 8'h56;
memory[16'h0c53] = 8'h5a;
memory[16'h0c54] = 8'h7f;
memory[16'h0c55] = 8'haf;
memory[16'h0c56] = 8'h70;
memory[16'h0c57] = 8'hfd;
memory[16'h0c58] = 8'h31;
memory[16'h0c59] = 8'h60;
memory[16'h0c5a] = 8'h0c;
memory[16'h0c5b] = 8'h7f;
memory[16'h0c5c] = 8'h1c;
memory[16'h0c5d] = 8'h0f;
memory[16'h0c5e] = 8'hc2;
memory[16'h0c5f] = 8'h20;
memory[16'h0c60] = 8'h56;
memory[16'h0c61] = 8'he2;
memory[16'h0c62] = 8'hf0;
memory[16'h0c63] = 8'heb;
memory[16'h0c64] = 8'h07;
memory[16'h0c65] = 8'h1a;
memory[16'h0c66] = 8'hf7;
memory[16'h0c67] = 8'h52;
memory[16'h0c68] = 8'hd0;
memory[16'h0c69] = 8'h50;
memory[16'h0c6a] = 8'hfd;
memory[16'h0c6b] = 8'haf;
memory[16'h0c6c] = 8'h42;
memory[16'h0c6d] = 8'hdd;
memory[16'h0c6e] = 8'heb;
memory[16'h0c6f] = 8'hf9;
memory[16'h0c70] = 8'hdc;
memory[16'h0c71] = 8'h80;
memory[16'h0c72] = 8'h3c;
memory[16'h0c73] = 8'h40;
memory[16'h0c74] = 8'h26;
memory[16'h0c75] = 8'he3;
memory[16'h0c76] = 8'h10;
memory[16'h0c77] = 8'h90;
memory[16'h0c78] = 8'he2;
memory[16'h0c79] = 8'hfb;
memory[16'h0c7a] = 8'hf9;
memory[16'h0c7b] = 8'h42;
memory[16'h0c7c] = 8'h13;
memory[16'h0c7d] = 8'h0c;
memory[16'h0c7e] = 8'h0f;
memory[16'h0c7f] = 8'hc2;
memory[16'h0c80] = 8'h30;
memory[16'h0c81] = 8'h0c;
memory[16'h0c82] = 8'hff;
memory[16'h0c83] = 8'h1c;
memory[16'h0c84] = 8'hff;
memory[16'h0c85] = 8'h82;
memory[16'h0c86] = 8'h20;
memory[16'h0c87] = 8'ha6;
memory[16'h0c88] = 8'he3;
memory[16'h0c89] = 8'h15;
memory[16'h0c8a] = 8'h6b;
memory[16'h0c8b] = 8'h12;
memory[16'h0c8c] = 8'h42;
memory[16'h0c8d] = 8'h22;
memory[16'h0c8e] = 8'heb;
memory[16'h0c8f] = 8'h0a;
memory[16'h0c90] = 8'hb6;
memory[16'h0c91] = 8'he3;
memory[16'h0c92] = 8'h10;
memory[16'h0c93] = 8'ha6;
memory[16'h0c94] = 8'he3;
memory[16'h0c95] = 8'h1d;
memory[16'h0c96] = 8'heb;
memory[16'h0c97] = 8'h02;
memory[16'h0c98] = 8'h3c;
memory[16'h0c99] = 8'h7f;
memory[16'h0c9a] = 8'h42;
memory[16'h0c9b] = 8'hd3;
memory[16'h0c9c] = 8'h2c;
memory[16'h0c9d] = 8'h00;
memory[16'h0c9e] = 8'h60;
memory[16'h0c9f] = 8'he2;
memory[16'h0ca0] = 8'h92;
memory[16'h0ca1] = 8'h20;
memory[16'h0ca2] = 8'h8b;
memory[16'h0ca3] = 8'hc5;
memory[16'h0ca4] = 8'h28;
memory[16'h0ca5] = 8'he0;
memory[16'h0ca6] = 8'h38;
memory[16'h0ca7] = 8'he1;
memory[16'h0ca8] = 8'h82;
memory[16'h0ca9] = 8'h72;
memory[16'h0caa] = 8'ha0;
memory[16'h0cab] = 8'he2;
memory[16'h0cac] = 8'h42;
memory[16'h0cad] = 8'h77;
memory[16'h0cae] = 8'heb;
memory[16'h0caf] = 8'hf8;
memory[16'h0cb0] = 8'h92;
memory[16'h0cb1] = 8'h72;
memory[16'h0cb2] = 8'h80;
memory[16'h0cb3] = 8'he2;
memory[16'h0cb4] = 8'ha2;
memory[16'h0cb5] = 8'h31;
memory[16'h0cb6] = 8'h6b;
memory[16'h0cb7] = 8'h08;
memory[16'h0cb8] = 8'h80;
memory[16'h0cb9] = 8'he2;
memory[16'h0cba] = 8'h82;
memory[16'h0cbb] = 8'h72;
memory[16'h0cbc] = 8'ha0;
memory[16'h0cbd] = 8'he2;
memory[16'h0cbe] = 8'h8b;
memory[16'h0cbf] = 8'hf0;
memory[16'h0cc0] = 8'ha2;
memory[16'h0cc1] = 8'h02;
memory[16'h0cc2] = 8'h7b;
memory[16'h0cc3] = 8'hf4;
memory[16'h0cc4] = 8'h92;
memory[16'h0cc5] = 8'h60;
memory[16'h0cc6] = 8'ha0;
memory[16'h0cc7] = 8'he0;
memory[16'h0cc8] = 8'haf;
memory[16'h0cc9] = 8'hd6;
memory[16'h0cca] = 8'h0c;
memory[16'h0ccb] = 8'ha4;
memory[16'h0ccc] = 8'h6b;
memory[16'h0ccd] = 8'h08;
memory[16'h0cce] = 8'hd6;
memory[16'h0ccf] = 8'h08;
memory[16'h0cd0] = 8'h24;
memory[16'h0cd1] = 8'h68;
memory[16'h0cd2] = 8'h5a;
memory[16'h0cd3] = 8'ha6;
memory[16'h0cd4] = 8'he6;
memory[16'h0cd5] = 8'h60;
memory[16'h0cd6] = 8'haf;
memory[16'h0cd7] = 8'hd6;
memory[16'h0cd8] = 8'h0c;
memory[16'h0cd9] = 8'hc9;
memory[16'h0cda] = 8'h6b;
memory[16'h0cdb] = 8'hfa;
memory[16'h0cdc] = 8'ha6;
memory[16'h0cdd] = 8'he6;
memory[16'h0cde] = 8'h20;
memory[16'h0cdf] = 8'heb;
memory[16'h0ce0] = 8'hf2;
memory[16'h0ce1] = 8'hd6;
memory[16'h0ce2] = 8'h0c;
memory[16'h0ce3] = 8'hce;
memory[16'h0ce4] = 8'h8b;
memory[16'h0ce5] = 8'hf6;
memory[16'h0ce6] = 8'ha0;
memory[16'h0ce7] = 8'he0;
memory[16'h0ce8] = 8'h82;
memory[16'h0ce9] = 8'h60;
memory[16'h0cea] = 8'h69;
memory[16'h0ceb] = 8'h5a;
memory[16'h0cec] = 8'hd6;
memory[16'h0ced] = 8'h08;
memory[16'h0cee] = 8'h27;
memory[16'h0cef] = 8'h42;
memory[16'h0cf0] = 8'h66;
memory[16'h0cf1] = 8'heb;
memory[16'h0cf2] = 8'he0;
memory[16'h0cf3] = 8'haf;
memory[16'h0cf4] = 8'hd6;
memory[16'h0cf5] = 8'h0d;
memory[16'h0cf6] = 8'h32;
memory[16'h0cf7] = 8'hfb;
memory[16'h0cf8] = 8'h71;
memory[16'h0cf9] = 8'hd6;
memory[16'h0cfa] = 8'h0d;
memory[16'h0cfb] = 8'h09;
memory[16'h0cfc] = 8'heb;
memory[16'h0cfd] = 8'h58;
memory[16'h0cfe] = 8'hd4;
memory[16'h0cff] = 8'h6e;
memory[16'h0d00] = 8'hfb;
memory[16'h0d01] = 8'h68;
memory[16'h0d02] = 8'hd6;
memory[16'h0d03] = 8'h0d;
memory[16'h0d04] = 8'h09;
memory[16'h0d05] = 8'h6b;
memory[16'h0d06] = 8'h2b;
memory[16'h0d07] = 8'h8b;
memory[16'h0d08] = 8'h2d;
memory[16'h0d09] = 8'ha6;
memory[16'h0d0a] = 8'he6;
memory[16'h0d0b] = 8'h3c;
memory[16'h0d0c] = 8'h6b;
memory[16'h0d0d] = 8'h5c;
memory[16'h0d0e] = 8'ha6;
memory[16'h0d0f] = 8'he6;
memory[16'h0d10] = 8'h3d;
memory[16'h0d11] = 8'h6b;
memory[16'h0d12] = 8'h57;
memory[16'h0d13] = 8'ha6;
memory[16'h0d14] = 8'he6;
memory[16'h0d15] = 8'h3e;
memory[16'h0d16] = 8'haf;
memory[16'h0d17] = 8'ha6;
memory[16'h0d18] = 8'h6f;
memory[16'h0d19] = 8'he6;
memory[16'h0d1a] = 8'h6b;
memory[16'h0d1b] = 8'h03;
memory[16'h0d1c] = 8'he6;
memory[16'h0d1d] = 8'h6f;
memory[16'h0d1e] = 8'hc9;
memory[16'h0d1f] = 8'hd4;
memory[16'h0d20] = 8'h6e;
memory[16'h0d21] = 8'hfb;
memory[16'h0d22] = 8'h47;
memory[16'h0d23] = 8'ha6;
memory[16'h0d24] = 8'he6;
memory[16'h0d25] = 8'h22;
memory[16'h0d26] = 8'heb;
memory[16'h0d27] = 8'hf7;
memory[16'h0d28] = 8'ha6;
memory[16'h0d29] = 8'h6f;
memory[16'h0d2a] = 8'he6;
memory[16'h0d2b] = 8'h6b;
memory[16'h0d2c] = 8'h03;
memory[16'h0d2d] = 8'he6;
memory[16'h0d2e] = 8'h6f;
memory[16'h0d2f] = 8'hd7;
memory[16'h0d30] = 8'h30;
memory[16'h0d31] = 8'h6e;
memory[16'h0d32] = 8'hd4;
memory[16'h0d33] = 8'h6e;
memory[16'h0d34] = 8'hfb;
memory[16'h0d35] = 8'h34;
memory[16'h0d36] = 8'hd6;
memory[16'h0d37] = 8'h0d;
memory[16'h0d38] = 8'h58;
memory[16'h0d39] = 8'hfb;
memory[16'h0d3a] = 8'h2f;
memory[16'h0d3b] = 8'hac;
memory[16'h0d3c] = 8'h03;
memory[16'h0d3d] = 8'hbc;
memory[16'h0d3e] = 8'hc1;
memory[16'h0d3f] = 8'hdc;
memory[16'h0d40] = 8'h03;
memory[16'h0d41] = 8'hd6;
memory[16'h0d42] = 8'h03;
memory[16'h0d43] = 8'haf;
memory[16'h0d44] = 8'h6b;
memory[16'h0d45] = 8'hec;
memory[16'h0d46] = 8'ha6;
memory[16'h0d47] = 8'he6;
memory[16'h0d48] = 8'h24;
memory[16'h0d49] = 8'heb;
memory[16'h0d4a] = 8'h1e;
memory[16'h0d4b] = 8'hd4;
memory[16'h0d4c] = 8'h6e;
memory[16'h0d4d] = 8'hfb;
memory[16'h0d4e] = 8'h1b;
memory[16'h0d4f] = 8'hdc;
memory[16'h0d50] = 8'h03;
memory[16'h0d51] = 8'hd6;
memory[16'h0d52] = 8'h03;
memory[16'h0d53] = 8'haf;
memory[16'h0d54] = 8'h6b;
memory[16'h0d55] = 8'hdc;
memory[16'h0d56] = 8'hcf;
memory[16'h0d57] = 8'haf;
memory[16'h0d58] = 8'ha6;
memory[16'h0d59] = 8'he6;
memory[16'h0d5a] = 8'h28;
memory[16'h0d5b] = 8'heb;
memory[16'h0d5c] = 8'h0e;
memory[16'h0d5d] = 8'hd6;
memory[16'h0d5e] = 8'h0d;
memory[16'h0d5f] = 8'h32;
memory[16'h0d60] = 8'hfb;
memory[16'h0d61] = 8'h08;
memory[16'h0d62] = 8'ha6;
memory[16'h0d63] = 8'he6;
memory[16'h0d64] = 8'h29;
memory[16'h0d65] = 8'heb;
memory[16'h0d66] = 8'hef;
memory[16'h0d67] = 8'h30;
memory[16'h0d68] = 8'h6e;
memory[16'h0d69] = 8'hdf;
memory[16'h0d6a] = 8'haf;
memory[16'h0d6b] = 8'hd6;
memory[16'h0d6c] = 8'h03;
memory[16'h0d6d] = 8'hd9;
memory[16'h0d6e] = 8'hfb;
memory[16'h0d6f] = 8'h1e;
memory[16'h0d70] = 8'hd4;
memory[16'h0d71] = 8'h6e;
memory[16'h0d72] = 8'hfb;
memory[16'h0d73] = 8'hf6;
memory[16'h0d74] = 8'hd6;
memory[16'h0d75] = 8'h03;
memory[16'h0d76] = 8'he2;
memory[16'h0d77] = 8'hfb;
memory[16'h0d78] = 8'hf0;
memory[16'h0d79] = 8'hd4;
memory[16'h0d7a] = 8'h6e;
memory[16'h0d7b] = 8'hfb;
memory[16'h0d7c] = 8'hed;
memory[16'h0d7d] = 8'ha6;
memory[16'h0d7e] = 8'he6;
memory[16'h0d7f] = 8'h3b;
memory[16'h0d80] = 8'h6b;
memory[16'h0d81] = 8'he7;
memory[16'h0d82] = 8'ha6;
memory[16'h0d83] = 8'he6;
memory[16'h0d84] = 8'h0d;
memory[16'h0d85] = 8'h6b;
memory[16'h0d86] = 8'he2;
memory[16'h0d87] = 8'ha6;
memory[16'h0d88] = 8'he6;
memory[16'h0d89] = 8'h5d;
memory[16'h0d8a] = 8'heb;
memory[16'h0d8b] = 8'hed;
memory[16'h0d8c] = 8'h30;
memory[16'h0d8d] = 8'h6e;
memory[16'h0d8e] = 8'h4c;
memory[16'h0d8f] = 8'h05;
memory[16'h0d90] = 8'hd6;
memory[16'h0d91] = 8'h03;
memory[16'h0d92] = 8'he7;
memory[16'h0d93] = 8'h7b;
memory[16'h0d94] = 8'h18;
memory[16'h0d95] = 8'ha6;
memory[16'h0d96] = 8'he6;
memory[16'h0d97] = 8'h2d;
memory[16'h0d98] = 8'h6b;
memory[16'h0d99] = 8'h12;
memory[16'h0d9a] = 8'ha6;
memory[16'h0d9b] = 8'he6;
memory[16'h0d9c] = 8'h25;
memory[16'h0d9d] = 8'heb;
memory[16'h0d9e] = 8'hb7;
memory[16'h0d9f] = 8'hd4;
memory[16'h0da0] = 8'h6e;
memory[16'h0da1] = 8'hfb;
memory[16'h0da2] = 8'hc7;
memory[16'h0da3] = 8'hd6;
memory[16'h0da4] = 8'h03;
memory[16'h0da5] = 8'hf2;
memory[16'h0da6] = 8'hfb;
memory[16'h0da7] = 8'h10;
memory[16'h0da8] = 8'h4a;
memory[16'h0da9] = 8'hf5;
memory[16'h0daa] = 8'hcf;
memory[16'h0dab] = 8'haf;
memory[16'h0dac] = 8'h4e;
memory[16'h0dad] = 8'hd4;
memory[16'h0dae] = 8'h6e;
memory[16'h0daf] = 8'hfb;
memory[16'h0db0] = 8'hb9;
memory[16'h0db1] = 8'hd6;
memory[16'h0db2] = 8'h03;
memory[16'h0db3] = 8'he7;
memory[16'h0db4] = 8'hfb;
memory[16'h0db5] = 8'h02;
memory[16'h0db6] = 8'h4a;
memory[16'h0db7] = 8'hf5;
memory[16'h0db8] = 8'hef;
memory[16'h0db9] = 8'haf;
memory[16'h0dba] = 8'h02;
memory[16'h0dbb] = 8'h27;
memory[16'h0dbc] = 8'h0d;
memory[16'h0dbd] = 8'h37;
memory[16'h0dbe] = 8'h23;
memory[16'h0dbf] = 8'h23;
memory[16'h0dc0] = 8'h0d;
memory[16'h0dc1] = 8'h0d;
memory[16'h0dc2] = 8'h27;
memory[16'h0dc3] = 8'h0d;
memory[16'h0dc4] = 8'h23;
memory[16'h0dc5] = 8'h23;
memory[16'h0dc6] = 8'h3a;
memory[16'h0dc7] = 8'h23;
memory[16'h0dc8] = 8'h60;
memory[16'h0dc9] = 8'h60;
memory[16'h0dca] = 8'h50;
memory[16'h0dcb] = 8'hff;
memory[16'h0dcc] = 8'he6;
memory[16'h0dcd] = 8'h5a;
memory[16'h0dce] = 8'h41;
memory[16'h0dcf] = 8'hd6;
memory[16'h0dd0] = 8'h0b;
memory[16'h0dd1] = 8'h95;
memory[16'h0dd2] = 8'hb0;
memory[16'h0dd3] = 8'h58;
memory[16'h0dd4] = 8'hd4;
memory[16'h0dd5] = 8'h6e;
memory[16'h0dd6] = 8'hfb;
memory[16'h0dd7] = 8'h13;
memory[16'h0dd8] = 8'h2c;
memory[16'h0dd9] = 8'h07;
memory[16'h0dda] = 8'h3c;
memory[16'h0ddb] = 8'hc8;
memory[16'h0ddc] = 8'hdc;
memory[16'h0ddd] = 8'h17;
memory[16'h0dde] = 8'hc3;
memory[16'h0ddf] = 8'hd2;
memory[16'h0de0] = 8'h20;
memory[16'h0de1] = 8'h58;
memory[16'h0de2] = 8'ha2;
memory[16'h0de3] = 8'h67;
memory[16'h0de4] = 8'h6b;
memory[16'h0de5] = 8'h06;
memory[16'h0de6] = 8'ha6;
memory[16'h0de7] = 8'h58;
memory[16'h0de8] = 8'h12;
memory[16'h0de9] = 8'h7b;
memory[16'h0dea] = 8'hf1;
memory[16'h0deb] = 8'haf;
memory[16'h0dec] = 8'h38;
memory[16'h0ded] = 8'h58;
memory[16'h0dee] = 8'h06;
memory[16'h0def] = 8'he3;
memory[16'h0df0] = 8'hb9;
memory[16'h0df1] = 8'he6;
memory[16'h0df2] = 8'h5c;
memory[16'h0df3] = 8'hff;
memory[16'h0df4] = 8'hd6;
memory[16'h0df5] = 8'h08;
memory[16'h0df6] = 8'h78;
memory[16'h0df7] = 8'hd6;
memory[16'h0df8] = 8'h0b;
memory[16'h0df9] = 8'hf2;
memory[16'h0dfa] = 8'h2c;
memory[16'h0dfb] = 8'h0d;
memory[16'h0dfc] = 8'h4c;
memory[16'h0dfd] = 8'h0e;
memory[16'h0dfe] = 8'hc2;
memory[16'h0dff] = 8'h52;
memory[16'h0e00] = 8'h30;
memory[16'h0e01] = 8'he4;
memory[16'h0e02] = 8'hd4;
memory[16'h0e03] = 8'h6e;
memory[16'h0e04] = 8'hd6;
memory[16'h0e05] = 8'h03;
memory[16'h0e06] = 8'hd9;
memory[16'h0e07] = 8'hfb;
memory[16'h0e08] = 8'he2;
memory[16'h0e09] = 8'hd4;
memory[16'h0e0a] = 8'h6e;
memory[16'h0e0b] = 8'h6c;
memory[16'h0e0c] = 8'h3d;
memory[16'h0e0d] = 8'hd6;
memory[16'h0e0e] = 8'h0d;
memory[16'h0e0f] = 8'h32;
memory[16'h0e10] = 8'hfb;
memory[16'h0e11] = 8'hd9;
memory[16'h0e12] = 8'ha6;
memory[16'h0e13] = 8'he6;
memory[16'h0e14] = 8'h2c;
memory[16'h0e15] = 8'h6b;
memory[16'h0e16] = 8'heb;
memory[16'h0e17] = 8'ha6;
memory[16'h0e18] = 8'he6;
memory[16'h0e19] = 8'h3b;
memory[16'h0e1a] = 8'h6b;
memory[16'h0e1b] = 8'hb0;
memory[16'h0e1c] = 8'ha6;
memory[16'h0e1d] = 8'he6;
memory[16'h0e1e] = 8'h0d;
memory[16'h0e1f] = 8'h6b;
memory[16'h0e20] = 8'h14;
memory[16'h0e21] = 8'hcf;
memory[16'h0e22] = 8'haf;
memory[16'h0e23] = 8'hd4;
memory[16'h0e24] = 8'h6e;
memory[16'h0e25] = 8'h8b;
memory[16'h0e26] = 8'hf0;
memory[16'h0e27] = 8'hd4;
memory[16'h0e28] = 8'h6e;
memory[16'h0e29] = 8'hfb;
memory[16'h0e2a] = 8'hc0;
memory[16'h0e2b] = 8'ha6;
memory[16'h0e2c] = 8'he6;
memory[16'h0e2d] = 8'h3b;
memory[16'h0e2e] = 8'h6b;
memory[16'h0e2f] = 8'h9c;
memory[16'h0e30] = 8'ha6;
memory[16'h0e31] = 8'he6;
memory[16'h0e32] = 8'h0d;
memory[16'h0e33] = 8'heb;
memory[16'h0e34] = 8'hf2;
memory[16'h0e35] = 8'hdf;
memory[16'h0e36] = 8'haf;
memory[16'h0e37] = 8'h5c;
memory[16'h0e38] = 8'h00;
memory[16'h0e39] = 8'h0d;
memory[16'h0e3a] = 8'h5c;
memory[16'h0e3b] = 8'h01;
memory[16'h0e3c] = 8'hd6;
memory[16'h0e3d] = 8'h0c;
memory[16'h0e3e] = 8'hf4;
memory[16'h0e3f] = 8'hfb;
memory[16'h0e40] = 8'haa;
memory[16'h0e41] = 8'h42;
memory[16'h0e42] = 8'h55;
memory[16'h0e43] = 8'heb;
memory[16'h0e44] = 8'hc8;
memory[16'h0e45] = 8'h6c;
memory[16'h0e46] = 8'h3b;
memory[16'h0e47] = 8'he6;
memory[16'h0e48] = 8'h58;
memory[16'h0e49] = 8'h13;
memory[16'h0e4a] = 8'hd6;
memory[16'h0e4b] = 8'h0b;
memory[16'h0e4c] = 8'hf2;
memory[16'h0e4d] = 8'h8d;
memory[16'h0e4e] = 8'h0d;
memory[16'h0e4f] = 8'hcc;
memory[16'h0e50] = 8'hd4;
memory[16'h0e51] = 8'h6e;
memory[16'h0e52] = 8'ha6;
memory[16'h0e53] = 8'he6;
memory[16'h0e54] = 8'h22;
memory[16'h0e55] = 8'heb;
memory[16'h0e56] = 8'h03;
memory[16'h0e57] = 8'hd6;
memory[16'h0e58] = 8'h0d;
memory[16'h0e59] = 8'h17;
memory[16'h0e5a] = 8'hd6;
memory[16'h0e5b] = 8'h03;
memory[16'h0e5c] = 8'hd9;
memory[16'h0e5d] = 8'h7b;
memory[16'h0e5e] = 8'hc4;
memory[16'h0e5f] = 8'haf;
memory[16'h0e60] = 8'hd4;
memory[16'h0e61] = 8'h6e;
memory[16'h0e62] = 8'ha6;
memory[16'h0e63] = 8'he6;
memory[16'h0e64] = 8'h22;
memory[16'h0e65] = 8'heb;
memory[16'h0e66] = 8'h03;
memory[16'h0e67] = 8'hd6;
memory[16'h0e68] = 8'h0d;
memory[16'h0e69] = 8'h17;
memory[16'h0e6a] = 8'ha6;
memory[16'h0e6b] = 8'he6;
memory[16'h0e6c] = 8'h3b;
memory[16'h0e6d] = 8'h6b;
memory[16'h0e6e] = 8'hde;
memory[16'h0e6f] = 8'ha6;
memory[16'h0e70] = 8'he6;
memory[16'h0e71] = 8'h0d;
memory[16'h0e72] = 8'h6b;
memory[16'h0e73] = 8'hc1;
memory[16'h0e74] = 8'hd6;
memory[16'h0e75] = 8'h0d;
memory[16'h0e76] = 8'h36;
memory[16'h0e77] = 8'hfb;
memory[16'h0e78] = 8'ha8;
memory[16'h0e79] = 8'ha6;
memory[16'h0e7a] = 8'he6;
memory[16'h0e7b] = 8'h2c;
memory[16'h0e7c] = 8'heb;
memory[16'h0e7d] = 8'h99;
memory[16'h0e7e] = 8'h8b;
memory[16'h0e7f] = 8'he0;
memory[16'h0e80] = 8'hd6;
memory[16'h0e81] = 8'h0a;
memory[16'h0e82] = 8'hd4;
memory[16'h0e83] = 8'he6;
memory[16'h0e84] = 8'h58;
memory[16'h0e85] = 8'h12;
memory[16'h0e86] = 8'hd6;
memory[16'h0e87] = 8'h0b;
memory[16'h0e88] = 8'hf2;
memory[16'h0e89] = 8'hb0;
memory[16'h0e8a] = 8'he2;
memory[16'h0e8b] = 8'h38;
memory[16'h0e8c] = 8'h0e;
memory[16'h0e8d] = 8'h56;
memory[16'h0e8e] = 8'he3;
memory[16'h0e8f] = 8'hf0;
memory[16'h0e90] = 8'hf0;
memory[16'h0e91] = 8'he3;
memory[16'h0e92] = 8'hd6;
memory[16'h0e93] = 8'h0a;
memory[16'h0e94] = 8'ha3;
memory[16'h0e95] = 8'h8d;
memory[16'h0e96] = 8'h0a;
memory[16'h0e97] = 8'hd4;
memory[16'h0e98] = 8'hcc;
memory[16'h0e99] = 8'h45;
memory[16'h0e9a] = 8'h54;
memory[16'h0e9b] = 8'hd0;
memory[16'h0e9c] = 8'h52;
memory[16'h0e9d] = 8'h4f;
memory[16'h0e9e] = 8'h43;
memory[16'h0e9f] = 8'hc7;
memory[16'h0ea0] = 8'h4f;
memory[16'h0ea1] = 8'h54;
memory[16'h0ea2] = 8'h4f;
memory[16'h0ea3] = 8'hc9;
memory[16'h0ea4] = 8'h46;
memory[16'h0ea5] = 8'hc5;
memory[16'h0ea6] = 8'h4c;
memory[16'h0ea7] = 8'h53;
memory[16'h0ea8] = 8'h45;
memory[16'h0ea9] = 8'hd2;
memory[16'h0eaa] = 8'h45;
memory[16'h0eab] = 8'h54;
memory[16'h0eac] = 8'h55;
memory[16'h0ead] = 8'h52;
memory[16'h0eae] = 8'h4e;
memory[16'h0eaf] = 8'hc7;
memory[16'h0eb0] = 8'h4f;
memory[16'h0eb1] = 8'h53;
memory[16'h0eb2] = 8'h55;
memory[16'h0eb3] = 8'h42;
memory[16'h0eb4] = 8'hd7;
memory[16'h0eb5] = 8'h41;
memory[16'h0eb6] = 8'h49;
memory[16'h0eb7] = 8'h54;
memory[16'h0eb8] = 8'hd2;
memory[16'h0eb9] = 8'h45;
memory[16'h0eba] = 8'h4d;
memory[16'h0ebb] = 8'hc3;
memory[16'h0ebc] = 8'h41;
memory[16'h0ebd] = 8'h4c;
memory[16'h0ebe] = 8'h4c;
memory[16'h0ebf] = 8'hd3;
memory[16'h0ec0] = 8'h54;
memory[16'h0ec1] = 8'h4f;
memory[16'h0ec2] = 8'h50;
memory[16'h0ec3] = 8'hc5;
memory[16'h0ec4] = 8'h4e;
memory[16'h0ec5] = 8'h44;
memory[16'h0ec6] = 8'hd4;
memory[16'h0ec7] = 8'h52;
memory[16'h0ec8] = 8'h41;
memory[16'h0ec9] = 8'h50;
memory[16'h0eca] = 8'hd4;
memory[16'h0ecb] = 8'h4f;
memory[16'h0ecc] = 8'h46;
memory[16'h0ecd] = 8'h46;
memory[16'h0ece] = 8'hd0;
memory[16'h0ecf] = 8'h52;
memory[16'h0ed0] = 8'h49;
memory[16'h0ed1] = 8'h4e;
memory[16'h0ed2] = 8'h54;
memory[16'h0ed3] = 8'hd0;
memory[16'h0ed4] = 8'h54;
memory[16'h0ed5] = 8'h48;
memory[16'h0ed6] = 8'hc9;
memory[16'h0ed7] = 8'h4e;
memory[16'h0ed8] = 8'h50;
memory[16'h0ed9] = 8'h55;
memory[16'h0eda] = 8'h54;
memory[16'h0edb] = 8'hc5;
memory[16'h0edc] = 8'h52;
memory[16'h0edd] = 8'h52;
memory[16'h0ede] = 8'h4f;
memory[16'h0edf] = 8'h52;
memory[16'h0ee0] = 8'h8b;
memory[16'h0ee1] = 8'h54;
memory[16'h0ee2] = 8'h48;
memory[16'h0ee3] = 8'h45;
memory[16'h0ee4] = 8'h4e;
memory[16'h0ee5] = 8'hc3;
memory[16'h0ee6] = 8'h4f;
memory[16'h0ee7] = 8'h4d;
memory[16'h0ee8] = 8'h50;
memory[16'h0ee9] = 8'h20;
memory[16'h0eea] = 8'h4a;
memory[16'h0eeb] = 8'h55;
memory[16'h0eec] = 8'h2b;
memory[16'h0eed] = 8'h54;
memory[16'h0eee] = 8'h45;
memory[16'h0eef] = 8'h20;
memory[16'h0ef0] = 8'h52;
memory[16'h0ef1] = 8'h20;
memory[16'h0ef2] = 8'h5c;
memory[16'h0ef3] = 8'h5c;
memory[16'h0ef4] = 8'h5c;
memory[16'h0ef5] = 8'h5c;
memory[16'h0ef6] = 8'h5c;
memory[16'h0ef7] = 8'h5c;
memory[16'h0ef8] = 8'h5c;
memory[16'h0ef9] = 8'h5c;
memory[16'h0efa] = 8'h5c;
memory[16'h0efb] = 8'h5c;
memory[16'h0efc] = 8'h5c;
memory[16'h0efd] = 8'h5c;
memory[16'h0efe] = 8'h0a;
memory[16'h0eff] = 8'hff;
memory[16'h0f00] = 8'h00;
memory[16'h0f01] = 8'h20;
memory[16'h0f02] = 8'h59;
memory[16'h0f03] = 8'h58;
memory[16'h0f04] = 8'h43;
memory[16'h0f05] = 8'h56;
memory[16'h0f06] = 8'h42;
memory[16'h0f07] = 8'h4e;
memory[16'h0f08] = 8'h4d;
memory[16'h0f09] = 8'h2c;
memory[16'h0f0a] = 8'h2e;
memory[16'h0f0b] = 8'h2f;
memory[16'h0f0c] = 8'h0d;
memory[16'h0f0d] = 8'h1b;
memory[16'h0f0e] = 8'h00;
memory[16'h0f0f] = 8'h00;
memory[16'h0f10] = 8'h00;
memory[16'h0f11] = 8'h15;
memory[16'h0f12] = 8'h41;
memory[16'h0f13] = 8'h53;
memory[16'h0f14] = 8'h44;
memory[16'h0f15] = 8'h46;
memory[16'h0f16] = 8'h47;
memory[16'h0f17] = 8'h48;
memory[16'h0f18] = 8'h4a;
memory[16'h0f19] = 8'h4b;
memory[16'h0f1a] = 8'h4c;
memory[16'h0f1b] = 8'h2a;
memory[16'h0f1c] = 8'h2d;
memory[16'h0f1d] = 8'h0a;
memory[16'h0f1e] = 8'h00;
memory[16'h0f1f] = 8'h00;
memory[16'h0f20] = 8'h00;
memory[16'h0f21] = 8'h0b;
memory[16'h0f22] = 8'h51;
memory[16'h0f23] = 8'h57;
memory[16'h0f24] = 8'h45;
memory[16'h0f25] = 8'h52;
memory[16'h0f26] = 8'h54;
memory[16'h0f27] = 8'h5a;
memory[16'h0f28] = 8'h55;
memory[16'h0f29] = 8'h49;
memory[16'h0f2a] = 8'h4f;
memory[16'h0f2b] = 8'h50;
memory[16'h0f2c] = 8'h2b;
memory[16'h0f2d] = 8'h0b;
memory[16'h0f2e] = 8'h00;
memory[16'h0f2f] = 8'h00;
memory[16'h0f30] = 8'h00;
memory[16'h0f31] = 8'h0a;
memory[16'h0f32] = 8'h31;
memory[16'h0f33] = 8'h32;
memory[16'h0f34] = 8'h33;
memory[16'h0f35] = 8'h34;
memory[16'h0f36] = 8'h35;
memory[16'h0f37] = 8'h36;
memory[16'h0f38] = 8'h37;
memory[16'h0f39] = 8'h38;
memory[16'h0f3a] = 8'h39;
memory[16'h0f3b] = 8'h30;
memory[16'h0f3c] = 8'h08;
memory[16'h0f3d] = 8'h1a;
memory[16'h0f3e] = 8'h00;
memory[16'h0f3f] = 8'h00;
memory[16'h0f40] = 8'hff;
memory[16'h0f41] = 8'hff;
memory[16'h0f42] = 8'hff;
memory[16'h0f43] = 8'hdd;
memory[16'h0f44] = 8'hdf;
memory[16'h0f45] = 8'hdf;
memory[16'h0f46] = 8'haa;
memory[16'h0f47] = 8'hff;
memory[16'h0f48] = 8'hff;
memory[16'h0f49] = 8'h50;
memory[16'h0f4a] = 8'h50;
memory[16'h0f4b] = 8'h5f;
memory[16'h0f4c] = 8'h69;
memory[16'h0f4d] = 8'h69;
memory[16'h0f4e] = 8'h6f;
memory[16'h0f4f] = 8'h6d;
memory[16'h0f50] = 8'hb7;
memory[16'h0f51] = 8'h6f;
memory[16'h0f52] = 8'h6d;
memory[16'h0f53] = 8'hb7;
memory[16'h0f54] = 8'haf;
memory[16'h0f55] = 8'hdd;
memory[16'h0f56] = 8'hff;
memory[16'h0f57] = 8'hff;
memory[16'h0f58] = 8'hdb;
memory[16'h0f59] = 8'hbb;
memory[16'h0f5a] = 8'hdf;
memory[16'h0f5b] = 8'hbd;
memory[16'h0f5c] = 8'hdd;
memory[16'h0f5d] = 8'hbf;
memory[16'h0f5e] = 8'h69;
memory[16'h0f5f] = 8'h09;
memory[16'h0f60] = 8'h6f;
memory[16'h0f61] = 8'hfd;
memory[16'h0f62] = 8'h8d;
memory[16'h0f63] = 8'hff;
memory[16'h0f64] = 8'hff;
memory[16'h0f65] = 8'hfd;
memory[16'h0f66] = 8'hbf;
memory[16'h0f67] = 8'hff;
memory[16'h0f68] = 8'h0f;
memory[16'h0f69] = 8'hff;
memory[16'h0f6a] = 8'hff;
memory[16'h0f6b] = 8'hff;
memory[16'h0f6c] = 8'hbf;
memory[16'h0f6d] = 8'hed;
memory[16'h0f6e] = 8'hb7;
memory[16'h0f6f] = 8'h7f;
memory[16'h0f70] = 8'h94;
memory[16'h0f71] = 8'h62;
memory[16'h0f72] = 8'h9f;
memory[16'h0f73] = 8'hd9;
memory[16'h0f74] = 8'hdd;
memory[16'h0f75] = 8'h8f;
memory[16'h0f76] = 8'h1e;
memory[16'h0f77] = 8'h97;
memory[16'h0f78] = 8'h0f;
memory[16'h0f79] = 8'h1e;
memory[16'h0f7a] = 8'h9e;
memory[16'h0f7b] = 8'h1f;
memory[16'h0f7c] = 8'h75;
memory[16'h0f7d] = 8'h0d;
memory[16'h0f7e] = 8'hdf;
memory[16'h0f7f] = 8'h07;
memory[16'h0f80] = 8'h1e;
memory[16'h0f81] = 8'h1f;
memory[16'h0f82] = 8'h97;
memory[16'h0f83] = 8'h16;
memory[16'h0f84] = 8'h9f;
memory[16'h0f85] = 8'h0e;
memory[16'h0f86] = 8'hdb;
memory[16'h0f87] = 8'hbf;
memory[16'h0f88] = 8'h96;
memory[16'h0f89] = 8'h96;
memory[16'h0f8a] = 8'h9f;
memory[16'h0f8b] = 8'h96;
memory[16'h0f8c] = 8'h8e;
memory[16'h0f8d] = 8'h9f;
memory[16'h0f8e] = 8'hfb;
memory[16'h0f8f] = 8'hfb;
memory[16'h0f90] = 8'hff;
memory[16'h0f91] = 8'hfd;
memory[16'h0f92] = 8'hfd;
memory[16'h0f93] = 8'hbf;
memory[16'h0f94] = 8'hdb;
memory[16'h0f95] = 8'h7b;
memory[16'h0f96] = 8'hdf;
memory[16'h0f97] = 8'hf0;
memory[16'h0f98] = 8'hf0;
memory[16'h0f99] = 8'hff;
memory[16'h0f9a] = 8'hbd;
memory[16'h0f9b] = 8'hed;
memory[16'h0f9c] = 8'hbf;
memory[16'h0f9d] = 8'h96;
memory[16'h0f9e] = 8'hdf;
memory[16'h0f9f] = 8'hdf;
memory[16'h0fa0] = 8'h86;
memory[16'h0fa1] = 8'h47;
memory[16'h0fa2] = 8'h8f;
memory[16'h0fa3] = 8'h96;
memory[16'h0fa4] = 8'h60;
memory[16'h0fa5] = 8'h6f;
memory[16'h0fa6] = 8'h16;
memory[16'h0fa7] = 8'h16;
memory[16'h0fa8] = 8'h1f;
memory[16'h0fa9] = 8'h87;
memory[16'h0faa] = 8'h77;
memory[16'h0fab] = 8'h8f;
memory[16'h0fac] = 8'h16;
memory[16'h0fad] = 8'h66;
memory[16'h0fae] = 8'h1f;
memory[16'h0faf] = 8'h07;
memory[16'h0fb0] = 8'h17;
memory[16'h0fb1] = 8'h0f;
memory[16'h0fb2] = 8'h07;
memory[16'h0fb3] = 8'h17;
memory[16'h0fb4] = 8'h7f;
memory[16'h0fb5] = 8'h87;
memory[16'h0fb6] = 8'h46;
memory[16'h0fb7] = 8'h8f;
memory[16'h0fb8] = 8'h66;
memory[16'h0fb9] = 8'h06;
memory[16'h0fba] = 8'h6f;
memory[16'h0fbb] = 8'h8d;
memory[16'h0fbc] = 8'hdd;
memory[16'h0fbd] = 8'h8f;
memory[16'h0fbe] = 8'h0e;
memory[16'h0fbf] = 8'he6;
memory[16'h0fc0] = 8'h9f;
memory[16'h0fc1] = 8'h65;
memory[16'h0fc2] = 8'h35;
memory[16'h0fc3] = 8'h6f;
memory[16'h0fc4] = 8'h77;
memory[16'h0fc5] = 8'h77;
memory[16'h0fc6] = 8'h0f;
memory[16'h0fc7] = 8'h60;
memory[16'h0fc8] = 8'h06;
memory[16'h0fc9] = 8'h6f;
memory[16'h0fca] = 8'h62;
memory[16'h0fcb] = 8'h46;
memory[16'h0fcc] = 8'h6f;
memory[16'h0fcd] = 8'h96;
memory[16'h0fce] = 8'h66;
memory[16'h0fcf] = 8'h9f;
memory[16'h0fd0] = 8'h16;
memory[16'h0fd1] = 8'h17;
memory[16'h0fd2] = 8'h7f;
memory[16'h0fd3] = 8'h96;
memory[16'h0fd4] = 8'h64;
memory[16'h0fd5] = 8'h8f;
memory[16'h0fd6] = 8'h16;
memory[16'h0fd7] = 8'h15;
memory[16'h0fd8] = 8'h6f;
memory[16'h0fd9] = 8'h87;
memory[16'h0fda] = 8'h9e;
memory[16'h0fdb] = 8'h1f;
memory[16'h0fdc] = 8'h8d;
memory[16'h0fdd] = 8'hdd;
memory[16'h0fde] = 8'hdf;
memory[16'h0fdf] = 8'h66;
memory[16'h0fe0] = 8'h66;
memory[16'h0fe1] = 8'h9f;
memory[16'h0fe2] = 8'haa;
memory[16'h0fe3] = 8'haa;
memory[16'h0fe4] = 8'hdf;
memory[16'h0fe5] = 8'h66;
memory[16'h0fe6] = 8'h00;
memory[16'h0fe7] = 8'h9f;
memory[16'h0fe8] = 8'h66;
memory[16'h0fe9] = 8'h96;
memory[16'h0fea] = 8'h6f;
memory[16'h0feb] = 8'haa;
memory[16'h0fec] = 8'hdd;
memory[16'h0fed] = 8'hdf;
memory[16'h0fee] = 8'h0d;
memory[16'h0fef] = 8'hb7;
memory[16'h0ff0] = 8'h0f;
memory[16'h0ff1] = 8'h9b;
memory[16'h0ff2] = 8'hbb;
memory[16'h0ff3] = 8'h9f;
memory[16'h0ff4] = 8'hf0;
memory[16'h0ff5] = 8'h66;
memory[16'h0ff6] = 8'h0f;
memory[16'h0ff7] = 8'h9d;
memory[16'h0ff8] = 8'hdd;
memory[16'h0ff9] = 8'h9f;
memory[16'h0ffa] = 8'h7b;
memory[16'h0ffb] = 8'hde;
memory[16'h0ffc] = 8'hef;
memory[16'h0ffd] = 8'hff;
memory[16'h0ffe] = 8'hff;
memory[16'h0fff] = 8'h0f;
