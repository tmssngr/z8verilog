initial begin
	if (isRom) begin
		`include "memory.vh"
	end
end
