    @(negedge clk);

#1000000
