localparam FETCH_MSB = 3;
localparam FETCH_INC  = 4'b1;
localparam FETCH_INSTR0  = 0;
localparam FETCH_INSTR1  = FETCH_INSTR0 + 1;
localparam FETCH_INSTR2  = FETCH_INSTR1 + 1;
localparam FETCH_SECOND0 = FETCH_INSTR2 + 1;
localparam FETCH_SECOND1 = FETCH_SECOND0 + 1;
localparam FETCH_SECOND2 = FETCH_SECOND1 + 1;
localparam FETCH_THIRD0  = FETCH_SECOND2 + 1;
localparam FETCH_THIRD1  = FETCH_THIRD0 + 1;
localparam FETCH_THIRD2  = FETCH_THIRD1 + 1;
localparam FETCH_DECODE  = FETCH_THIRD2 + 1;

localparam OP_MSB = 4;
localparam OP_UNDECIDED = 0;
localparam OP_DECODE    = OP_UNDECIDED + 1;
localparam OP_LD        = OP_DECODE + 1;
localparam OP_ALU1      = OP_LD + 1;
localparam OP_ALU1DA    = OP_ALU1 + 1;
localparam OP_ALU1WORD  = OP_ALU1DA + 1;
localparam OP_ALU2      = OP_ALU1WORD + 1;
localparam OP_POP       = OP_ALU2 + 1;
localparam OP_PUSH      = OP_POP + 1;
localparam OP_DJNZ      = OP_PUSH + 1;
localparam OP_JP        = OP_DJNZ + 1;
localparam OP_JR        = OP_JP + 1;
localparam OP_JP_IRR    = OP_JR + 1;
localparam OP_CALL      = OP_JP_IRR + 1;
localparam OP_RET       = OP_CALL + 1;
localparam OP_IRET      = OP_RET + 1;
localparam OP_LDC       = OP_IRET + 1;
localparam OP_MISC      = OP_LDC + 1;
localparam OP_ISR       = OP_MISC + 1;
localparam OP_ILLEGAL   = OP_ISR + 1;

localparam OPSTATE_MSB = 3;
localparam OPSTATE_INC = 4'b1;
localparam OPSTATE0 = 0;
localparam OPSTATE1 = OPSTATE0 + 1;
localparam OPSTATE2 = OPSTATE1 + 1;
localparam OPSTATE3 = OPSTATE2 + 1;
localparam OPSTATE4 = OPSTATE3 + 1;
localparam OPSTATE5 = OPSTATE4 + 1;
localparam OPSTATE6 = OPSTATE5 + 1;
localparam OPSTATE7 = OPSTATE6 + 1;
localparam OPSTATE8 = OPSTATE7 + 1;
localparam OPSTATE9 = OPSTATE8 + 1;
localparam OPSTATE10 = OPSTATE9 + 1;

localparam SIO_IDLE  = 0;
localparam SIO_START = SIO_IDLE  + 1;
localparam SIO_BIT0  = SIO_START + 1;
localparam SIO_BIT1  = SIO_BIT0  + 1;
localparam SIO_BIT2  = SIO_BIT1  + 1;
localparam SIO_BIT3  = SIO_BIT2  + 1;
localparam SIO_BIT4  = SIO_BIT3  + 1;
localparam SIO_BIT5  = SIO_BIT4  + 1;
localparam SIO_BIT6  = SIO_BIT5  + 1;
localparam SIO_BIT7  = SIO_BIT6  + 1;
localparam SIO_STOP1 = SIO_BIT7  + 1;
localparam SIO_STOP2 = SIO_STOP1 + 1;
