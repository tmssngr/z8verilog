localparam FLAG_INDEX_C = 7;
localparam FLAG_INDEX_Z = 6;
localparam FLAG_INDEX_S = 5;
localparam FLAG_INDEX_V = 4;
localparam FLAG_INDEX_D = 3; // 1 after sub, 0 after add
localparam FLAG_INDEX_H = 2; // half-carry
